----------------------------------------------------------------------------------------------------------------------------------------------------------------
-- LSD.TOS, April 2017 (DO NOT REMOVE THIS LINE)
--
-- Blop sound ROM (dual port, synchronous read). At 48kHz, this sound has a duration of about 85 miliseconds.
--
-- The blop sound was kindly put in the public domain by Mark DiAngelo (http://soundbible.com/2067-Blop.html).
--
-- Octave/matlab commands used to generate the data for the ROM:
--   x=wavread('Blop-Mark_DiAngelo-79054334.wav'); % read the .wav file
--   i=2496;                                       % index of the first sample we are interested in
--   y=round(65536*x(i:i+4095,1));                 % convert 4096 samples to integers (in this case, in the range -32767 to 32767)
--   y(end)=0;                                     % make sure the last sample is zero (silence)
--   save blop.txt y                               % save y
-- The 16-bit integers stored in the file blop.txt were then converted to hexadecimal and, after that, to VHDL.
--

library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

entity blop_sound_rom is
  port
  (
    clock : in std_logic;

    addr0_0 : in  std_logic_vector(11 downto 0); -- sample number
    data0_1 : out std_logic_vector(15 downto 0); -- sample value (available with a delay of one clock cycle)

    addr1_0 : in  std_logic_vector(11 downto 0); -- sample number
    data1_1 : out std_logic_vector(15 downto 0)  -- sample value (available with a delay of one clock cycle)
  );
end blop_sound_rom;

architecture v1 of blop_sound_rom is
  --
  -- The sound samples (to be interpreted as 16-bit signed integers)
  --
  type rom_t is array(0 to 4095) of std_logic_vector(15 downto 0);
  constant sound_data : rom_t :=
  (
    x"0004",x"0005",x"FFFE",x"FFFF",x"0009",x"0003",x"FFFC",x"FFF8",x"FFF7",x"FFF9",x"0001",x"0002",x"FFFF",x"FFFD",x"FFFE",x"FFF5",
    x"FFF2",x"FFF5",x"FFFD",x"FFF5",x"FFFE",x"FFFE",x"FFF8",x"FFF8",x"FFF6",x"FFEF",x"FFF7",x"FFFC",x"FFFE",x"FFFB",x"FFFA",x"FFF4",
    x"FFE8",x"FFE6",x"FFEB",x"FFF7",x"FFFD",x"0002",x"0003",x"FFF6",x"FFEF",x"FFE9",x"FFE8",x"FFEB",x"FFED",x"FFEC",x"FFE7",x"FFF0",
    x"FFF7",x"FFEF",x"FFE9",x"FFE1",x"FFDE",x"FFE7",x"FFE8",x"FFEA",x"FFE7",x"FFED",x"FFE9",x"FFEB",x"FFE5",x"FFDC",x"FFDE",x"FFDE",
    x"FFE2",x"FFD5",x"FFDA",x"FFD3",x"FFD7",x"FFD6",x"FFD7",x"FFCF",x"FFC1",x"FFBE",x"FFC3",x"FFCA",x"FFCE",x"FFCA",x"FFB7",x"FFB4",
    x"FFC0",x"FFD4",x"FFCE",x"FFCC",x"FFB9",x"FFB2",x"FFB4",x"FFB6",x"FFB5",x"FFC3",x"FFBF",x"FFB3",x"FFC1",x"FFC4",x"FFC9",x"FFCF",
    x"FFC2",x"FFAF",x"FF9F",x"FFAC",x"FFB6",x"FFAA",x"FFB2",x"FFBB",x"FFB9",x"FFB8",x"FFB0",x"FFAC",x"FFA0",x"FFB0",x"FFC6",x"FFBE",
    x"FFC1",x"FFB3",x"FF96",x"FF96",x"FFB6",x"FFC7",x"FFCB",x"FFC0",x"FFA3",x"FF7E",x"FF7E",x"FF8C",x"FFAB",x"FFC5",x"FFC4",x"FFC0",
    x"FFC2",x"FF97",x"FF91",x"FFA7",x"FFAC",x"FFCB",x"FFD8",x"FFC5",x"FFB6",x"FFC5",x"FFC5",x"FFC8",x"FFD4",x"FFD1",x"FFC5",x"FFB9",
    x"FFB3",x"FFC2",x"FFCC",x"FFD5",x"FFDB",x"FFD1",x"FFD9",x"FFCC",x"FFCE",x"FFD6",x"FFEB",x"FFFD",x"000D",x"FFF9",x"FFF3",x"FFD5",
    x"FFEA",x"FFF2",x"FFF4",x"001D",x"0003",x"0002",x"FFFC",x"0000",x"000C",x"0005",x"0012",x"0021",x"004C",x"0067",x"005C",x"003C",
    x"001A",x"0013",x"0025",x"0042",x"003C",x"0040",x"005B",x"001C",x"000A",x"0002",x"0017",x"0006",x"0002",x"0029",x"001E",x"FFB7",
    x"FF65",x"FF4E",x"FF26",x"FEE8",x"FE97",x"FE0A",x"FD2A",x"FC43",x"FB22",x"FA13",x"F8C2",x"F75C",x"F5BB",x"F40A",x"F275",x"F061",
    x"EE60",x"EC68",x"EA72",x"E832",x"E555",x"E0F9",x"DB79",x"D684",x"D398",x"D343",x"D46A",x"D45F",x"D2FF",x"D073",x"CDDE",x"CC0C",
    x"CB8C",x"CBF7",x"CC29",x"CC63",x"CCD1",x"CC87",x"CB95",x"CB34",x"CB2C",x"CAF1",x"CB93",x"CD24",x"CE6D",x"CE69",x"CDF0",x"CFA0",
    x"D1A8",x"D2F0",x"D4EC",x"D643",x"D7E2",x"D97E",x"DC02",x"DFDC",x"E074",x"E0E9",x"E3E7",x"E8E7",x"ECF1",x"EFC0",x"F231",x"F663",
    x"FA01",x"FEF1",x"0461",x"0934",x"0E34",x"13CC",x"1A29",x"1FF7",x"258B",x"29CA",x"2E63",x"33B8",x"38C1",x"3F1A",x"4466",x"48EF",
    x"4D4D",x"5219",x"56E1",x"5AF3",x"5F71",x"63AA",x"685B",x"6D93",x"70A6",x"736C",x"7588",x"766D",x"7795",x"7761",x"75B1",x"736C",
    x"704C",x"6C04",x"666C",x"5F81",x"57F0",x"4F63",x"4651",x"3C8B",x"3219",x"26E6",x"1B6E",x"102C",x"050D",x"F850",x"EBAE",x"E050",
    x"D471",x"C8BA",x"BDA7",x"B30A",x"A9A5",x"A258",x"9C23",x"9645",x"9286",x"9034",x"902B",x"922A",x"95D1",x"9A00",x"A02A",x"A7DA",
    x"B032",x"B995",x"C3E5",x"CE6D",x"DA00",x"E633",x"F28B",x"FF56",x"0C0C",x"18F6",x"25F4",x"32A2",x"3E28",x"4901",x"53AB",x"5D2D",
    x"65F7",x"6D2C",x"72A7",x"7601",x"7771",x"770E",x"750F",x"71AC",x"6C21",x"655C",x"5DCC",x"5482",x"4A12",x"3EB3",x"3268",x"25A4",
    x"18D2",x"0B13",x"FC79",x"EEB8",x"E1DD",x"D4E3",x"C861",x"BC6B",x"B16C",x"A851",x"A0D0",x"9A5C",x"95E9",x"936A",x"9296",x"9419",
    x"9739",x"9B06",x"A062",x"A790",x"B03F",x"B987",x"C367",x"CE23",x"D9CB",x"E611",x"F2AD",x"FF15",x"0B57",x"17AF",x"2410",x"3016",
    x"3B0A",x"454A",x"4EC6",x"56B9",x"5CF0",x"61D1",x"64D1",x"65E1",x"6580",x"638C",x"5FE8",x"5A74",x"5389",x"4B5C",x"425E",x"3884",
    x"2D6F",x"2160",x"14E8",x"086A",x"FC24",x"EFA5",x"E301",x"D6C1",x"CB25",x"C03E",x"B626",x"AD84",x"A6B4",x"A190",x"9E14",x"9C2E",
    x"9BD0",x"9D19",x"A016",x"A4B7",x"AADD",x"B21A",x"BA20",x"C396",x"CE5E",x"D975",x"E4C8",x"F090",x"FCB5",x"08BB",x"14D6",x"20D7",
    x"2C56",x"3748",x"41BC",x"4B2C",x"530B",x"5994",x"5ECB",x"6269",x"6449",x"6487",x"62F4",x"5FB7",x"5B11",x"553E",x"4DCF",x"44A9",
    x"3A8C",x"2FF2",x"2497",x"1874",x"0BFC",x"FF44",x"F28D",x"E621",x"D9D6",x"CDE7",x"C2CF",x"B8D4",x"B024",x"A8E7",x"A32D",x"9EFE",
    x"9C52",x"9B50",x"9C3C",x"9EC6",x"A2CD",x"A810",x"AEC2",x"B6F2",x"C018",x"C9CC",x"D41C",x"DF3F",x"EB0F",x"F73A",x"0327",x"0F0B",
    x"1AFC",x"267D",x"3154",x"3B51",x"4461",x"4C60",x"5324",x"585C",x"5BF5",x"5DFD",x"5E81",x"5D8B",x"5AFC",x"56EA",x"5139",x"4A10",
    x"41C3",x"3896",x"2E96",x"23C6",x"184C",x"0C5F",x"0048",x"F430",x"E846",x"DC84",x"D136",x"C688",x"BD11",x"B534",x"AED0",x"A981",
    x"A55B",x"A2C8",x"A232",x"A343",x"A5A3",x"A94E",x"AE64",x"B4D4",x"BC7D",x"C50D",x"CEA5",x"D8EA",x"E385",x"EE88",x"F9C2",x"053F",
    x"10EF",x"1C69",x"2749",x"3161",x"3ACB",x"4340",x"4A67",x"5055",x"551A",x"5863",x"59FF",x"5A45",x"5928",x"5649",x"51AC",x"4BD5",
    x"4503",x"3D12",x"33F7",x"29F0",x"1F5A",x"148D",x"0958",x"FDAC",x"F18B",x"E5AC",x"DA9D",x"D056",x"C6DF",x"BE44",x"B6A6",x"B053",
    x"AB5D",x"A7F0",x"A5D4",x"A542",x"A66F",x"A94E",x"AD9F",x"B2B7",x"B8BB",x"C004",x"C861",x"D190",x"DB41",x"E57D",x"F05D",x"FB61",
    x"0635",x"10E8",x"1B51",x"254A",x"2E9F",x"3707",x"3E59",x"44C8",x"4A4C",x"4E87",x"50FF",x"5203",x"51B0",x"4FDC",x"4CB7",x"486A",
    x"42FB",x"3C77",x"34E9",x"2C5F",x"2329",x"1952",x"0EFB",x"046E",x"F9D8",x"EF57",x"E531",x"DB8B",x"D29D",x"CAA7",x"C382",x"BD39",
    x"B830",x"B490",x"B276",x"B1BA",x"B23C",x"B40A",x"B6FF",x"BB2D",x"C049",x"C697",x"CE11",x"D653",x"DEF7",x"E7DA",x"F144",x"FB3A",
    x"051F",x"0EC3",x"1814",x"213C",x"2A00",x"31D6",x"38B3",x"3E83",x"430A",x"469F",x"4910",x"4A24",x"49DC",x"4859",x"45AB",x"419F",
    x"3C80",x"3671",x"2F91",x"27A7",x"1EDD",x"158C",x"0BD9",x"021E",x"F87B",x"EEEB",x"E550",x"DC0F",x"D391",x"CBF3",x"C547",x"BFA6",
    x"BB2F",x"B7E4",x"B5C3",x"B505",x"B59F",x"B77B",x"BA77",x"BE85",x"C38B",x"C95C",x"D025",x"D7DE",x"E03C",x"E8E3",x"F1E3",x"FB31",
    x"0482",x"0DCA",x"16E5",x"1FA0",x"27BB",x"2F1B",x"35C4",x"3B77",x"401B",x"439C",x"4604",x"470F",x"46CA",x"4587",x"4318",x"3F54",
    x"3A7A",x"34CC",x"2E3F",x"26BE",x"1EB7",x"162B",x"0D0E",x"039B",x"FA54",x"F14A",x"E885",x"DFE5",x"D7D9",x"D092",x"CA18",x"C49D",
    x"C067",x"BD49",x"BB47",x"BA77",x"BACC",x"BC4B",x"BEF9",x"C2BF",x"C780",x"CD07",x"D35B",x"DA65",x"E239",x"EA76",x"F314",x"FBDA",
    x"0480",x"0D1B",x"158A",x"1DB5",x"2548",x"2C27",x"3253",x"3792",x"3BC4",x"3EF8",x"412B",x"4226",x"41F2",x"408B",x"3E2C",x"3AC2",
    x"364B",x"30F1",x"2AAC",x"239C",x"1BEA",x"13D0",x"0B4B",x"029E",x"F9CD",x"F112",x"E890",x"E069",x"D8DB",x"D1F7",x"CBEF",x"C6CB",
    x"C2AD",x"BFAF",x"BDB9",x"BCD9",x"BD1C",x"BE89",x"C101",x"C453",x"C8A8",x"CDE0",x"D3D6",x"DA85",x"E1E4",x"E9AC",x"F1BB",x"FA05",
    x"025D",x"0AA6",x"12B6",x"1A7E",x"21D0",x"287A",x"2E77",x"339F",x"37F2",x"3B3B",x"3D6B",x"3EAC",x"3ED6",x"3DE0",x"3BF5",x"38FD",
    x"3506",x"302C",x"2A82",x"243B",x"1D49",x"15EC",x"0E1F",x"063E",x"FE2E",x"F62B",x"EE50",x"E6DB",x"DFBA",x"D958",x"D3B3",x"CED2",
    x"CAE2",x"C7D3",x"C5C9",x"C4CC",x"C4D0",x"C5D7",x"C7DC",x"CAB5",x"CE64",x"D2FF",x"D84B",x"DE27",x"E496",x"EB78",x"F292",x"F9DF",
    x"014C",x"08A4",x"0FC5",x"16A6",x"1D28",x"22FD",x"2827",x"2C9A",x"3050",x"332D",x"3508",x"360C",x"3629",x"3533",x"3343",x"309C",
    x"2D2B",x"28E8",x"23F8",x"1E62",x"183C",x"11BB",x"0AFB",x"0419",x"FD2E",x"F63F",x"EFA7",x"E95A",x"E380",x"DE1E",x"D99C",x"D5C8",
    x"D2B1",x"D07C",x"CF37",x"CEC9",x"CF39",x"D099",x"D2DB",x"D5C6",x"D971",x"DDCB",x"E2C6",x"E832",x"EE14",x"F454",x"FABF",x"013A",
    x"07A7",x"0E04",x"142C",x"19ED",x"1F46",x"240E",x"2822",x"2B88",x"2E2F",x"2FF4",x"30E6",x"30E6",x"301A",x"2E67",x"2BD9",x"2883",
    x"247A",x"1FDA",x"1A87",x"14B5",x"0E7D",x"0817",x"0179",x"FABF",x"F40D",x"ED8B",x"E756",x"E178",x"DC23",x"D77D",x"D381",x"D03B",
    x"CDCC",x"CC34",x"CB6D",x"CB9C",x"CC99",x"CE74",x"D122",x"D4A2",x"D8BE",x"DD6B",x"E2B7",x"E887",x"EE9D",x"F4FC",x"FB99",x"0233",
    x"08BB",x"0F21",x"1552",x"1B17",x"2053",x"2510",x"2929",x"2C85",x"2F1B",x"3103",x"320E",x"324F",x"31AE",x"3040",x"2DFE",x"2AFB",
    x"2745",x"22FD",x"1E11",x"18A8",x"12D5",x"0CB9",x"0660",x"0012",x"F9BB",x"F3A5",x"EDBA",x"E83B",x"E327",x"DEB0",x"DAD3",x"D7A1",
    x"D530",x"D378",x"D284",x"D260",x"D2F4",x"D442",x"D648",x"D90C",x"DC6B",x"E055",x"E4BC",x"E99D",x"EED7",x"F440",x"F9DD",x"FF8B",
    x"0533",x"0AA3",x"0FEB",x"14E4",x"1966",x"1D72",x"20E9",x"23C6",x"25F7",x"277F",x"2854",x"2875",x"27E6",x"2691",x"24AF",x"2211",
    x"1ED6",x"1B22",x"1709",x"126E",x"0DAD",x"08AD",x"0371",x"FE40",x"F91A",x"F427",x"EF6F",x"EB08",x"E713",x"E3A4",x"E0D0",x"DE89",
    x"DCED",x"DBF6",x"DB94",x"DBDC",x"DCD4",x"DE63",x"E094",x"E35C",x"E69E",x"EA4C",x"EE77",x"F2E0",x"F782",x"FC55",x"0135",x"0623",
    x"0AE7",x"0F72",x"13BC",x"17B8",x"1B46",x"1E42",x"20DA",x"22D2",x"2419",x"24CD",x"24FC",x"2473",x"2339",x"2174",x"1F1C",x"1C41",
    x"18E4",x"1513",x"10ED",x"0C7E",x"07D8",x"0317",x"FE30",x"F964",x"F4A9",x"F037",x"EBFE",x"E829",x"E4D7",x"E1EF",x"DF8D",x"DDC6",
    x"DC9C",x"DC04",x"DC16",x"DCBC",x"DDF3",x"DFBF",x"E211",x"E4D1",x"E810",x"EBB2",x"EFA5",x"F3E4",x"F852",x"FCD7",x"0162",x"05F2",
    x"0A55",x"0E89",x"1280",x"160C",x"1939",x"1BEC",x"1E21",x"1FD1",x"20FB",x"217B",x"2180",x"20EE",x"1FC1",x"1E18",x"1BE5",x"1935",
    x"1619",x"129D",x"0EC7",x"0AC7",x"0696",x"0242",x"FDEF",x"F9B2",x"F587",x"F199",x"EE06",x"EAAA",x"E7CF",x"E56D",x"E389",x"E237",
    x"E154",x"E0FB",x"E135",x"E215",x"E368",x"E526",x"E74B",x"E9EB",x"ECF9",x"F068",x"F40F",x"F7E7",x"FBE7",x"FFFE",x"03FC",x"07FC",
    x"0BC7",x"0F67",x"12B4",x"15A2",x"1833",x"1A52",x"1BF0",x"1D0B",x"1DA8",x"1DB5",x"1D3E",x"1C48",x"1ADA",x"18EF",x"168C",x"13C1",
    x"10B0",x"0D56",x"09B3",x"05E9",x"01FD",x"FDFF",x"FA0A",x"F638",x"F272",x"EEFD",x"EBE4",x"E914",x"E6B5",x"E4C3",x"E361",x"E261",
    x"E1F8",x"E20E",x"E2A9",x"E3B6",x"E545",x"E73B",x"E99B",x"EC61",x"EF69",x"F2CA",x"F658",x"FA01",x"FDC7",x"019F",x"0565",x"090B",
    x"0C8E",x"0FDB",x"12E9",x"1599",x"17DE",x"19BB",x"1B10",x"1BFE",x"1C70",x"1C60",x"1BD3",x"1AC6",x"1952",x"1779",x"1535",x"1296",
    x"0FB3",x"0C8E",x"0938",x"05BA",x"022E",x"FEA0",x"FB1D",x"F7C3",x"F491",x"F189",x"EEC9",x"EC5F",x"EA62",x"E8D1",x"E7B0",x"E701",
    x"E6D0",x"E703",x"E7A9",x"E8C6",x"EA43",x"EC29",x"EE6B",x"F0E6",x"F39C",x"F67E",x"F98E",x"FCD5",x"0019",x"0349",x"066D",x"0979",
    x"0C52",x"0EF4",x"114F",x"1357",x"14FD",x"164B",x"1724",x"1792",x"1796",x"1731",x"1646",x"14FD",x"1350",x"1156",x"0F0D",x"0C75",
    x"09A6",x"06B5",x"0395",x"007B",x"FD57",x"FA2B",x"F716",x"F442",x"F19B",x"EF47",x"ED32",x"EB6F",x"EA16",x"E91F",x"E894",x"E875",
    x"E8C6",x"E982",x"EA9A",x"EC15",x"EDE5",x"F013",x"F275",x"F50E",x"F7E2",x"FACD",x"FDCB",x"00E5",x"03E8",x"06E2",x"09BC",x"0C71",
    x"0EF9",x"1139",x"1328",x"14B9",x"15F5",x"16D6",x"1755",x"1769",x"1710",x"1651",x"1537",x"13AF",x"11EE",x"0FC5",x"0D68",x"0ADE",
    x"0815",x"053A",x"0233",x"FF32",x"FC3C",x"F942",x"F677",x"F3DB",x"F17A",x"EF4B",x"ED8B",x"EC07",x"EAED",x"EA2C",x"E9C5",x"E9D7",
    x"EA3E",x"EB0A",x"EC30",x"EDAF",x"EF7D",x"F189",x"F3D4",x"F65A",x"F906",x"FBCE",x"FEAE",x"0184",x"045C",x"0720",x"09BF",x"0C30",
    x"0E6C",x"1066",x"121D",x"1379",x"1484",x"1530",x"1571",x"155B",x"14FD",x"142E",x"130F",x"1197",x"0FD2",x"0DDA",x"0BB9",x"094A",
    x"06C5",x"0422",x"0188",x"FEDA",x"FC47",x"F9BB",x"F757",x"F529",x"F32F",x"F185",x"F029",x"EF11",x"EE4E",x"EDDC",x"EDC1",x"EE06",
    x"EEAC",x"EFA5",x"F0F1",x"F275",x"F439",x"F634",x"F86D",x"FAB8",x"FD2A",x"FF97",x"0225",x"049B",x"06FD",x"0938",x"0B57",x"0D44",
    x"0EF2",x"105B",x"117A",x"123B",x"12C6",x"12FB",x"12DA",x"126E",x"11B0",x"1097",x"0F33",x"0D8B",x"0BAE",x"09A2",x"0766",x"051B",
    x"02B2",x"003F",x"FDBB",x"FB58",x"F90A",x"F6DA",x"F4DB",x"F311",x"F183",x"F03E",x"EF40",x"EE82",x"EE2A",x"EE26",x"EE6B",x"EEF2",
    x"EFD4",x"F101",x"F263",x"F411",x"F5E3",x"F7D9",x"F9FC",x"FC38",x"FE7A",x"00D9",x"0325",x"0565",x"0785",x"097E",x"0B47",x"0CE1",
    x"0E4C",x"0F6D",x"1047",x"10D2",x"1107",x"10EF",x"108A",x"0FE0",x"0EFB",x"0DC3",x"0C5B",x"0AB5",x"08DC",x"06D7",x"04B8",x"0288",
    x"003D",x"FE05",x"FBDC",x"F9BB",x"F7B1",x"F5CF",x"F421",x"F2C1",x"F180",x"F097",x"EFE6",x"EF7F",x"EF6D",x"EF9A",x"F020",x"F0EF",
    x"F1F3",x"F341",x"F4C0",x"F66C",x"F850",x"FA44",x"FC6B",x"FE9E",x"00D5",x"02F8",x"0502",x"06EF",x"08D8",x"0A91",x"0C13",x"0D58",
    x"0E60",x"0F35",x"0FB5",x"0FDD",x"0FC5",x"0F6D",x"0ED9",x"0DF3",x"0CCB",x"0B76",x"09DC",x"0817",x"062E",x"0419",x"01F6",x"FFCF",
    x"FDB7",x"FB9D",x"F98E",x"F7A6",x"F5D6",x"F439",x"F2D7",x"F1B2",x"F0DD",x"F03B",x"EFDD",x"EFC2",x"F003",x"F07F",x"F142",x"F23F",
    x"F37F",x"F4DF",x"F687",x"F859",x"FA42",x"FC41",x"FE5B",x"0077",x"0295",x"04A2",x"06A1",x"088C",x"0A4E",x"0BC4",x"0D0E",x"0E26",
    x"0EFF",x"0F96",x"0FEF",x"0FEF",x"0FC2",x"0F47",x"0E84",x"0D94",x"0C5F",x"0AFB",x"096C",x"07BD",x"05DE",x"03F1",x"01FF",x"FFF7",
    x"FDF8",x"FC0B",x"FA32",x"F864",x"F6D1",x"F568",x"F435",x"F338",x"F267",x"F209",x"F1CA",x"F1D3",x"F214",x"F2A8",x"F36D",x"F46F",
    x"F5A4",x"F70D",x"F8AC",x"FA61",x"FC38",x"FE17",x"000B",x"01F6",x"03D8",x"05AA",x"076F",x"0919",x"0A8B",x"0BD4",x"0CF5",x"0DD1",
    x"0E80",x"0EE0",x"0F04",x"0EE5",x"0E7D",x"0DE3",x"0D09",x"0BFA",x"0AB5",x"0946",x"07B4",x"05F0",x"0434",x"0252",x"0060",x"FE81",
    x"FCAA",x"FAE5",x"F935",x"F7A1",x"F634",x"F503",x"F401",x"F33E",x"F2C5",x"F277",x"F279",x"F2AA",x"F323",x"F3D7",x"F4B7",x"F5D4",
    x"F714",x"F884",x"FA0E",x"FBB8",x"FD78",x"FF3B",x"0106",x"02D4",x"0496",x"064C",x"07D4",x"093D",x"0A94",x"0BBE",x"0CA9",x"0D5A",
    x"0DDA",x"0E07",x"0E14",x"0DD5",x"0D61",x"0CB4",x"0BC7",x"0A9D",x"0943",x"07CD",x"0633",x"0487",x"02C2",x"00EE",x"FF2B",x"FD60",
    x"FB9B",x"F9E4",x"F855",x"F6EE",x"F5B2",x"F49C",x"F3B1",x"F30F",x"F29F",x"F272",x"F279",x"F2B6",x"F338",x"F3E6",x"F4D2",x"F5F1",
    x"F736",x"F893",x"FA13",x"FBBC",x"FD6F",x"FF30",x"00F4",x"02AE",x"0451",x"05E2",x"075B",x"08BD",x"09EB",x"0AEB",x"0BBE",x"0C64",
    x"0CD4",x"0D07",x"0D00",x"0CBB",x"0C37",x"0B91",x"0AB7",x"099F",x"0868",x"06FA",x"0589",x"03F1",x"023E",x"008D",x"FEDD",x"FD28",
    x"FB7E",x"F9EA",x"F86D",x"F724",x"F5F7",x"F4F1",x"F421",x"F37D",x"F311",x"F2D9",x"F302",x"F338",x"F3C0",x"F46D",x"F54B",x"F656",
    x"F780",x"F8C7",x"FA32",x"FBC1",x"FD5B",x"FEFE",x"00A1",x"0240",x"03D8",x"0567",x"06C7",x"0815",x"093A",x"0A41",x"0B08",x"0BA7",
    x"0C0C",x"0C42",x"0C40",x"0C01",x"0BAA",x"0B13",x"0A50",x"095E",x"0844",x"0718",x"05CA",x"0453",x"02CF",x"0157",x"FFE5",x"FE64",
    x"FCE7",x"FB7E",x"FA2B",x"F8F6",x"F7E0",x"F6EC",x"F62B",x"F595",x"F539",x"F517",x"F513",x"F549",x"F5A7",x"F632",x"F6F0",x"F7DC",
    x"F8D9",x"F9FE",x"FB3D",x"FC7D",x"FDDF",x"FF53",x"00BC",x"0230",x"038A",x"04DC",x"0623",x"073E",x"0842",x"092B",x"09DA",x"0A70",
    x"0AD5",x"0B04",x"0B1A",x"0AFF",x"0AAA",x"0A4A",x"09AF",x"08EA",x"0805",x"0708",x"05F6",x"04D1",x"0395",x"0250",x"010D",x"FFC8",
    x"FE95",x"FD60",x"FC45",x"FB2D",x"FA4D",x"F978",x"F8C9",x"F849",x"F7E7",x"F7BE",x"F7BA",x"F7BC",x"F804",x"F862",x"F8E8",x"F98E",
    x"FA48",x"FB26",x"FC16",x"FD23",x"FE2C",x"FF4D",x"0069",x"0182",x"0297",x"039B",x"0489",x"0569",x"062A",x"06C9",x"0754",x"07BD",
    x"0801",x"0827",x"0822",x"0801",x"07AE",x"073E",x"06AA",x"060D",x"0551",x"0479",x"0395",x"0297",x"019F",x"009F",x"FF9B",x"FE8E",
    x"FD9C",x"FCBC",x"FBDC",x"FB22",x"FA80",x"F9F3",x"F97A",x"F932",x"F90C",x"F91A",x"F932",x"F962",x"F9A7",x"FA20",x"FA9E",x"FB3F",
    x"FBFB",x"FCC3",x"FD95",x"FE76",x"FF58",x"0048",x"012F",x"0218",x"02F3",x"03C8",x"046E",x"0524",x"05B3",x"0623",x"067F",x"06BC",
    x"06DF",x"06E4",x"06C0",x"0681",x"062C",x"05BC",x"0531",x"049F",x"03F3",x"0340",x"026F",x"019C",x"00BA",x"FFDE",x"FEFA",x"FE20",
    x"FD50",x"FC79",x"FBC1",x"FB17",x"FA8C",x"FA19",x"F9B9",x"F978",x"F95D",x"F954",x"F96A",x"F97A",x"F9BB",x"FA19",x"FA8C",x"FAFE",
    x"FB8D",x"FC28",x"FCCC",x"FD7D",x"FE35",x"FEEA",x"FFA4",x"0063",x"0111",x"01B1",x"0237",x"02B9",x"0329",x"0395",x"03D8",x"0409",
    x"042D",x"0438",x"0432",x"0417",x"03E5",x"03B0",x"0363",x"030E",x"02B7",x"024B",x"01D9",x"015E",x"00E0",x"006C",x"FFFE",x"FF8E",
    x"FF2D",x"FED8",x"FE87",x"FE3D",x"FE0C",x"FDDF",x"FDBB",x"FDC2",x"FDCB",x"FDF6",x"FE2C",x"FE66",x"FEB0",x"FF12",x"FF75",x"FFE3",
    x"0043",x"00B8",x"0126",x"018F",x"01F8",x"024B",x"0297",x"02E6",x"0322",x"0349",x"0366",x"036F",x"0366",x"0351",x"033D",x"0303",
    x"02D2",x"027A",x"021C",x"01AE",x"0138",x"00B8",x"002F",x"FFB4",x"FF2D",x"FEB4",x"FE40",x"FDD2",x"FD6D",x"FD11",x"FCB7",x"FC82",
    x"FC50",x"FC38",x"FC31",x"FC33",x"FC4A",x"FC7B",x"FCBA",x"FD11",x"FD7F",x"FDFA",x"FE73",x"FEFA",x"FF8E",x"0026",x"00BC",x"0159",
    x"01EF",x"0281",x"030A",x"0387",x"0400",x"0458",x"04B4",x"04EE",x"0524",x"053C",x"053F",x"0524",x"04FB",x"04B6",x"0480",x"0412",
    x"0399",x"030E",x"0286",x"01F8",x"0147",x"009F",x"FFF9",x"FF56",x"FEC6",x"FE1A",x"FD8A",x"FD13",x"FC91",x"FC31",x"FBE3",x"FBA6",
    x"FB80",x"FB75",x"FB75",x"FB96",x"FBCE",x"FC0D",x"FC62",x"FCD0",x"FD50",x"FDE4",x"FE7C",x"FF20",x"FFD8",x"0082",x"0126",x"01CE",
    x"026B",x"0305",x"0397",x"0419",x"0485",x"04CA",x"0516",x"0538",x"0551",x"054C",x"052D",x"04EE",x"049B",x"0438",x"03C6",x"033D",
    x"02A3",x"0208",x"0157",x"0098",x"FFDC",x"FF19",x"FE68",x"FDB0",x"FCFD",x"FC59",x"FBCC",x"FB46",x"FAD6",x"FA73",x"FA27",x"FA01",
    x"F9DB",x"F9E4",x"FA05",x"FA34",x"FA7C",x"FAE1",x"FB65",x"FBE0",x"FC79",x"FD31",x"FDFA",x"FEAB",x"FF5F",x"001B",x"00D7",x"019A",
    x"0252",x"02FF",x"0395",x"041D",x"049F",x"0504",x"0560",x"059A",x"05D3",x"05E2",x"05CE",x"05A8",x"056E",x"0524",x"04BF",x"0444",
    x"03B6",x"0320",x"0278",x"01C9",x"011D",x"005E",x"FFA4",x"FEF5",x"FE58",x"FDB3",x"FD1C",x"FC94",x"FC21",x"FBC5",x"FB67",x"FB3D",
    x"FB12",x"FB07",x"FB12",x"FB2F",x"FB6A",x"FBA8",x"FC06",x"FC76",x"FCF2",x"FD8A",x"FE13",x"FE99",x"FF32",x"FFC6",x"005E",x"00EB",
    x"0172",x"01F8",x"0262",x"02C9",x"0329",x"0366",x"039E",x"03C6",x"03D6",x"03DA",x"03CD",x"03A4",x"037E",x"0334",x"02D4",x"0278",
    x"0208",x"019A",x"011F",x"0096",x"0024",x"FFA2",x"FF27",x"FEB0",x"FE3B",x"FDDB",x"FD88",x"FD40",x"FD06",x"FCDB",x"FCC0",x"FCB7",
    x"FCBC",x"FCD5",x"FCFF",x"FD35",x"FD78",x"FDD2",x"FE2C",x"FE8C",x"FF0C",x"FF8B",x"0009",x"007B",x"00F2",x"016B",x"01D9",x"024B",
    x"02A3",x"02E4",x"032E",x"0358",x"0373",x"0387",x"0387",x"037C",x"0363",x"0329",x"02E8",x"0295",x"0242",x"01DD",x"0176",x"0102",
    x"0082",x"0009",x"FF90",x"FF19",x"FEAB",x"FE35",x"FDC9",x"FD66",x"FD18",x"FCDE",x"FC9F",x"FC79",x"FC69",x"FC5E",x"FC7B",x"FC86",
    x"FCBA",x"FCED",x"FD31",x"FD88",x"FDEF",x"FE5D",x"FEBF",x"FF27",x"FFB4",x"0031",x"00A1",x"011D",x"0179",x"01D2",x"022C",x"026B",
    x"02A7",x"02D6",x"0305",x"030E",x"0310",x"0301",x"02E1",x"02B2",x"0278",x"0235",x"01E9",x"0182",x"011D",x"00B6",x"004C",x"FFE3",
    x"FF68",x"FF05",x"FEA9",x"FE42",x"FDF4",x"FDA5",x"FD57",x"FD25",x"FCF4",x"FCDB",x"FCCE",x"FCCE",x"FCE9",x"FD0F",x"FD45",x"FD88",
    x"FDD9",x"FE32",x"FE8E",x"FEF3",x"FF6E",x"FFE7",x"0067",x"00E5",x"0164",x"01D7",x"0254",x"02B7",x"0310",x"035F",x"0395",x"03CF",
    x"03FC",x"0405",x"0409",x"0403",x"03DF",x"03A7",x"0363",x"0313",x"02BB",x"024B",x"01D0",x"0162",x"00D3",x"0045",x"FFBD",x"FF41",
    x"FEB2",x"FE30",x"FDAE",x"FD3C",x"FCDE",x"FC79",x"FC33",x"FBF0",x"FBC5",x"FBAD",x"FBA4",x"FBAF",x"FBC8",x"FBF7",x"FC38",x"FC82",
    x"FCD7",x"FD3E",x"FDB3",x"FE2E",x"FEB0",x"FF2B",x"FFBD",x"0045",x"00E2",x"016D",x"01FD",x"026D",x"02DF",x"0340",x"038E",x"03D3",
    x"0409",x"0419",x"0426",x"0419",x"0410",x"03E1",x"03AB",x"036C",x"0322",x"02D6",x"025F",x"01F6",x"017F",x"0100",x"0084",x"0000",
    x"FF82",x"FF05",x"FE90",x"FE20",x"FDB7",x"FD64",x"FD16",x"FCDE",x"FC9F",x"FC7D",x"FC74",x"FC67",x"FC7D",x"FC98",x"FCBE",x"FCFB",
    x"FD47",x"FD9E",x"FDFF",x"FE6A",x"FED4",x"FF51",x"FFC1",x"002B",x"00A1",x"0114",x"016D",x"01C9",x"0213",x"025D",x"0297",x"02BB",
    x"02CF",x"02ED",x"02EA",x"02DF",x"02C0",x"0293",x"0256",x"0208",x"01B3",x"0160",x"00F2",x"0080",x"0019",x"FFAD",x"FF36",x"FEBF",
    x"FE4B",x"FDE4",x"FD8F",x"FD35",x"FCE9",x"FCB3",x"FC7F",x"FC5E",x"FC47",x"FC45",x"FC55",x"FC70",x"FCA6",x"FCE2",x"FD1C",x"FD6D",
    x"FDC2",x"FE27",x"FE8C",x"FF00",x"FF77",x"FFEE",x"0063",x"00E0",x"0160",x"01C3",x"0225",x"027F",x"02DD",x"031C",x"0346",x"0373",
    x"037C",x"0387",x"0381",x"0371",x"0349",x"0327",x"02E6",x"02A7",x"0262",x"0208",x"01A5",x"0145",x"00DE",x"0069",x"0007",x"FF99",
    x"FF30",x"FECF",x"FE7A",x"FE29",x"FDDB",x"FDAE",x"FD7A",x"FD62",x"FD52",x"FD57",x"FD6D",x"FD8F",x"FDA7",x"FDDF",x"FE20",x"FE52",
    x"FE99",x"FEF3",x"FF46",x"FFB2",x"0009",x"0069",x"00D0",x"011D",x"0174",x"01D0",x"020F",x"024B",x"028A",x"02AC",x"02C7",x"02CD",
    x"02D2",x"02BE",x"02B0",x"027A",x"0242",x"0201",x"01BE",x"0164",x"0116",x"00BF",x"0067",x"FFFC",x"FF9D",x"FF39",x"FEDA",x"FE81",
    x"FE2C",x"FDDD",x"FD9C",x"FD66",x"FD45",x"FD2C",x"FD28",x"FD28",x"FD31",x"FD47",x"FD6F",x"FD9E",x"FDE4",x"FE23",x"FE64",x"FEBB",
    x"FF12",x"FF68",x"FFD3",x"0024",x"0084",x"00D3",x"0118",x"016B",x"01B7",x"01E4",x"021A",x"023E",x"0252",x"025F",x"025F",x"0256",
    x"0237",x"0211",x"01DB",x"019A",x"0149",x"0100",x"00AA",x"0048",x"FFE5",x"FF7E",x"FF1E",x"FEC4",x"FE61",x"FE0C",x"FDB3",x"FD64",
    x"FD1F",x"FCF0",x"FCCC",x"FCB1",x"FCA3",x"FCAA",x"FCAF",x"FCC5",x"FCF6",x"FD28",x"FD62",x"FDB7",x"FE11",x"FE76",x"FEE3",x"FF48",
    x"FFB4",x"0024",x"0092",x"00FB",x"0160",x"01C5",x"021A",x"0281",x"02C0",x"02F1",x"0329",x"0342",x"0349",x"034D",x"0337",x"030A",
    x"02CB",x"027D",x"0237",x"01E6",x"0176",x"00FD",x"008B",x"0010",x"FF8E",x"FF07",x"FE87",x"FE0A",x"FD9E",x"FD2C",x"FCC5",x"FC70",
    x"FC12",x"FBCC",x"FBA8",x"FB80",x"FB77",x"FB79",x"FB99",x"FBBA",x"FBF7",x"FC4C",x"FC9F",x"FCF8",x"FD74",x"FDF6",x"FE87",x"FF22",
    x"FFB6",x"004A",x"00E0",x"0176",x"0206",x"0288",x"030C",x"037E",x"03EE",x"044D",x"0485",x"04A6",x"04C6",x"04CA",x"04BA",x"0492",
    x"0463",x"0410",x"03B0",x"034D",x"02D8",x"0259",x"01C5",x"0131",x"0094",x"000B",x"FF68",x"FED8",x"FE4F",x"FDD9",x"FD59",x"FCE0",
    x"FC70",x"FC1B",x"FBD1",x"FBA4",x"FB75",x"FB70",x"FB79",x"FB87",x"FBB1",x"FBF7",x"FC43",x"FC9D",x"FCF8",x"FD78",x"FDF4",x"FE81",
    x"FF0C",x"FFA6",x"0036",x"00BC",x"014E",x"01CE",x"0247",x"02B2",x"0322",x"036F",x"03BD",x"03F7",x"0412",x"0429",x"0424",x"0419",
    x"0403",x"03D1",x"038C",x"0337",x"02CF",x"0266",x"01F4",x"017F",x"00F9",x"0075",x"FFE7",x"FF65",x"FEE1",x"FE64",x"FDF1",x"FD8A",
    x"FD2C",x"FCD7",x"FC9D",x"FC55",x"FC3A",x"FC2D",x"FC35",x"FC3C",x"FC60",x"FC9F",x"FCE9",x"FD3C",x"FDAA",x"FE15",x"FE8E",x"FF03",
    x"FF82",x"0007",x"008B",x"010B",x"0176",x"01E9",x"023E",x"02A7",x"0303",x"0349",x"038E",x"03B0",x"03B6",x"03BB",x"039E",x"037C",
    x"034B",x"0301",x"02B5",x"0247",x"01D2",x"0157",x"00E7",x"005C",x"FFD5",x"FF4D",x"FEB9",x"FE37",x"FDC0",x"FD50",x"FCEB",x"FC86",
    x"FC47",x"FC00",x"FBCE",x"FBA8",x"FBB1",x"FBB1",x"FBCA",x"FBF7",x"FC2D",x"FC74",x"FCE2",x"FD47",x"FDC4",x"FE56",x"FED6",x"FF61",
    x"FFF7",x"008F",x"0123",x"01B5",x"023E",x"02B7",x"0325",x"0399",x"03F3",x"0434",x"046A",x"0485",x"049D",x"04AB",x"049B",x"0479",
    x"043D",x"03F3",x"0392",x"0329",x"02B2",x"0237",x"01BA",x"0116",x"0084",x"FFE7",x"FF4F",x"FEC2",x"FE2E",x"FDB0",x"FD31",x"FCC9",
    x"FC62",x"FC0F",x"FBBA",x"FB96",x"FB75",x"FB6C",x"FB7B",x"FB99",x"FBCE",x"FC0B",x"FC5E",x"FCCC",x"FD39",x"FDC0",x"FE4B",x"FEE6",
    x"FF7A",x"001F",x"00CE",x"015E",x"01F8",x"0286",x"0305",x"038A",x"03F5",x"0453",x"04A4",x"04E0",x"0518",x"052A",x"0524",x"0509",
    x"04E7",x"04A8",x"045C",x"0405",x"0381",x"0303",x"0288",x"01F2",x"015B",x"00B1",x"000B",x"FF58",x"FEC6",x"FE27",x"FD86",x"FD04",
    x"FC76",x"FC06",x"FBA6",x"FB53",x"FB20",x"FB02",x"FAEC",x"FAEA",x"FB02",x"FB31",x"FB72",x"FBBC",x"FC1F",x"FC9A",x"FD0F",x"FD91",
    x"FE15",x"FEB0",x"FF48",x"FFE1",x"0077",x"011D",x"01A3",x"022A",x"02B9",x"0330",x"03A2",x"03EC",x"043F",x"0470",x"0499",x"04B4",
    x"04BD",x"04AD",x"0489",x"045A",x"0419",x"03CB",x"036C",x"0310",x"02A5",x"0223",x"01B3",x"011D",x"0094",x"0000",x"FF73",x"FEFC",
    x"FE76",x"FE03",x"FD95",x"FD28",x"FCC9",x"FC86",x"FC55",x"FC31",x"FC18",x"FC0B",x"FC16",x"FC28",x"FC47",x"FC84",x"FCC9",x"FD13",
    x"FD54",x"FDAC",x"FE1A",x"FE83",x"FEF3",x"FF56",x"FFC8",x"0026",x"0096",x"00F7",x"015E",x"01AA",x"01FF",x"023E",x"0271",x"0297",
    x"02B2",x"02BE",x"02B9",x"02A5",x"028A",x"0268",x"0223",x"01F2",x"019C",x"015B",x"010F",x"00BF",x"006C",x"000D",x"FFB8",x"FF5F",
    x"FF12",x"FEBD",x"FE71",x"FE32",x"FDFC",x"FDC2",x"FDA5",x"FD8A",x"FD76",x"FD76",x"FD7A",x"FD93",x"FDAC",x"FDE4",x"FE11",x"FE3B",
    x"FE87",x"FECD",x"FF1E",x"FF6A",x"FFBB",x"0010",x"005E",x"00A4",x"0104",x"0143",x"0198",x"01D2",x"0206",x"022C",x"0256",x"0266",
    x"0283",x"0288",x"028A",x"028C",x"026D",x"0249",x"0215",x"01E0",x"019F",x"0155",x"0114",x"00C5",x"0072",x"001B",x"FFD1",x"FF7E",
    x"FF29",x"FEEF",x"FEA9",x"FE6F",x"FE3B",x"FE15",x"FE08",x"FDE6",x"FDDD",x"FDE2",x"FDF6",x"FDFA",x"FE1E",x"FE3D",x"FE5F",x"FE8A",
    x"FEBD",x"FEFA",x"FF34",x"FF73",x"FFCA",x"0014",x"005A",x"00AD",x"0106",x"015B",x"01A5",x"01CE",x"0208",x"0230",x"0259",x"0274",
    x"0281",x"0283",x"027D",x"0268",x"024B",x"022C",x"01FD",x"01D4",x"019F",x"0164",x"0126",x"00E2",x"0092",x"0045",x"FFFC",x"FFAD",
    x"FF5F",x"FF03",x"FEB4",x"FE71",x"FE35",x"FE08",x"FDCB",x"FDA7",x"FD8A",x"FD7A",x"FD7D",x"FD7A",x"FD7F",x"FD9C",x"FDBE",x"FDD6",
    x"FDF6",x"FE1C",x"FE58",x"FE8A",x"FEBD",x"FF00",x"FF3B",x"FF7C",x"FFC6",x"0009",x"004C",x"0086",x"00C7",x"00F7",x"012F",x"0152",
    x"0169",x"017F",x"0193",x"01A8",x"01AA",x"01A8",x"01A8",x"019A",x"0179",x"0170",x"0155",x"0135",x"0114",x"00F9",x"00D0",x"009F",
    x"0077",x"004C",x"0014",x"FFF7",x"FFC3",x"FF9D",x"FF85",x"FF71",x"FF51",x"FF3B",x"FF22",x"FF15",x"FF12",x"FF05",x"FF17",x"FF1B",
    x"FF29",x"FF30",x"FF46",x"FF5F",x"FF7A",x"FF90",x"FFA6",x"FFC8",x"FFF5",x"0012",x"0036",x"004C",x"0069",x"0086",x"0092",x"00A6",
    x"00C1",x"00B3",x"00A1",x"00A6",x"009B",x"0096",x"0089",x"0080",x"0063",x"0055",x"0043",x"002D",x"002B",x"0024",x"001B",x"FFFE",
    x"FFEE",x"FFCF",x"FFD3",x"FFBF",x"FFAD",x"FFA9",x"FF99",x"FF97",x"FF8E",x"FF90",x"FF99",x"FF92",x"FF99",x"FFA9",x"FFBB",x"FFC3",
    x"FFD8",x"FFE5",x"000B",x"001F",x"003A",x"0057",x"0063",x"006E",x"0098",x"00A4",x"00BA",x"00C5",x"00C7",x"00E5",x"00F2",x"00F9",
    x"00FD",x"00FD",x"010D",x"0102",x"0102",x"0100",x"00F0",x"00D5",x"00C1",x"00A6",x"0092",x"0089",x"0065",x"0055",x"002D",x"001B",
    x"0000",x"FFEE",x"FFCF",x"FFBF",x"FFA9",x"FF94",x"FF85",x"FF73",x"FF68",x"FF51",x"FF5A",x"FF5A",x"FF5C",x"FF5F",x"FF5F",x"FF68",
    x"FF73",x"FF90",x"FFA2",x"FFB8",x"FFD1",x"FFEC",x"0004",x"001D",x"003F",x"005C",x"007B",x"00A1",x"00B3",x"00D7",x"00EB",x"0108",
    x"0114",x"012F",x"0150",x"0157",x"0164",x"016D",x"0170",x"0174",x"016D",x"016B",x"0150",x"0149",x"0145",x"0133",x"0123",x"010B",
    x"00F9",x"00D9",x"00B6",x"0098",x"0080",x"005E",x"0041",x"0028",x"0007",x"FFF5",x"FFD8",x"FFC3",x"FFA6",x"FF9D",x"FF97",x"FF92",
    x"FF99",x"FF9B",x"FF95",x"FF9B",x"FFA0",x"FFB0",x"FFB2",x"FFBE",x"FFD8",x"FFF1",x"000D",x"000F",x"001A",x"0032",x"004E",x"0056",
    x"005D",x"006A",x"0079",x"0077",x"0080",x"0086",x"008E",x"0082",x"0077",x"006F",x"0061",x"004A",x"0040",x"0024",x"0014",x"FFF0",
    x"FFD2",x"FFB5",x"FF93",x"FF81",x"FF62",x"FF4F",x"FF2E",x"FF13",x"FEF0",x"FED5",x"FEBE",x"FEB4",x"FE98",x"FE93",x"FE95",x"FE8F",
    x"FE93",x"FE92",x"FE98",x"FEB0",x"FEC2",x"FED2",x"FEED",x"FF0A",x"FF1E",x"FF43",x"FF6B",x"FF8E",x"FFC0",x"FFE9",x"0017",x"0041",
    x"0077",x"00A5",x"00DB",x"010E",x"0138",x"0156",x"017C",x"019F",x"01C3",x"01C9",x"01D5",x"01EC",x"01F8",x"01F0",x"01E4",x"01DC",
    x"01CC",x"01BB",x"019A",x"0187",x"0163",x"0136",x"0111",x"00E2",x"00AF",x"0071",x"003A",x"0010",x"FFDE",x"FFA5",x"FF77",x"FF4E",
    x"FF1C",x"FEFF",x"FEDF",x"FEC1",x"FEAA",x"FE99",x"FE84",x"FE7A",x"FE72",x"FE76",x"FE79",x"FE7F",x"FE7C",x"FE99",x"FEA7",x"FEB7",
    x"FED4",x"FEFC",x"FF19",x"FF3F",x"FF71",x"FFA4",x"FFC4",x"FFEE",x"001B",x"0042",x"0071",x"0092",x"00B7",x"00D0",x"00F3",x"0109",
    x"0121",x"0127",x"0136",x"013B",x"0142",x"013D",x"0138",x"0134",x"011B",x"00FF",x"00E9",x"00D3",x"00B3",x"0090",x"0077",x"0056",
    x"0035",x"0015",x"FFF6",x"FFD9",x"FFB9",x"FF9D",x"FF80",x"FF6C",x"FF4F",x"FF44",x"FF33",x"FF26",x"FF23",x"FF24",x"FF26",x"FF2D",
    x"FF36",x"FF44",x"FF4D",x"FF5A",x"FF74",x"FF88",x"FFA3",x"FFBD",x"FFDB",x"FFF5",x"0012",x"0031",x"0048",x"0062",x"0070",x"0081",
    x"009D",x"00A8",x"00B8",x"00C2",x"00C8",x"00C5",x"00CB",x"00C7",x"00BF",x"00B9",x"00B4",x"00A3",x"0094",x"007D",x"0066",x"004C",
    x"0038",x"001F",x"0007",x"FFF3",x"FFD9",x"FFC4",x"FFAB",x"FF97",x"FF8A",x"FF76",x"FF76",x"FF65",x"FF5B",x"FF58",x"FF55",x"FF52",
    x"FF56",x"FF5D",x"FF65",x"FF72",x"FF81",x"FF92",x"FFA6",x"FFBD",x"FFD5",x"FFE7",x"0005",x"001C",x"0034",x"0048",x"005E",x"0076",
    x"0088",x"0098",x"00AD",x"00B6",x"00C1",x"00C6",x"00C6",x"00C9",x"00C3",x"00BB",x"00AF",x"009E",x"0092",x"007B",x"006A",x"0057",
    x"0043",x"0029",x"0013",x"FFFE",x"FFEB",x"FFD1",x"FFB8",x"FFA6",x"FF8D",x"FF7D",x"FF6D",x"FF60",x"FF55",x"FF50",x"FF4B",x"FF4A",
    x"FF48",x"FF4F",x"FF51",x"FF5A",x"FF67",x"FF78",x"FF86",x"FF99",x"FFAD",x"FFC5",x"FFDA",x"FFF5",x"000D",x"0022",x"0036",x"004D",
    x"0062",x"0073",x"0081",x"0092",x"00A0",x"00A7",x"00B4",x"00BC",x"00BE",x"00B9",x"00B5",x"00B5",x"00AB",x"00A2",x"0094",x"0088",
    x"0078",x"0064",x"004F",x"003F",x"002A",x"0014",x"FFFE",x"FFED",x"FFD5",x"FFBD",x"FFAE",x"FF9B",x"FF88",x"FF7C",x"FF71",x"FF66",
    x"FF5F",x"FF5C",x"FF59",x"FF5A",x"FF5E",x"FF68",x"FF6E",x"FF7A",x"FF87",x"FF95",x"FFA7",x"FFB7",x"FFC7",x"FFDD",x"FFEF",x"0001",
    x"0014",x"0027",x"0038",x"0045",x"0057",x"0063",x"006E",x"0078",x"0081",x"0084",x"0089",x"008D",x"008E",x"0088",x"0085",x"0080",
    x"0075",x"0068",x"005C",x"004D",x"0043",x"0031",x"001E",x"0015",x"0002",x"FFF4",x"FFE9",x"FFD9",x"FFCD",x"FFC0",x"FFBA",x"FFB4",
    x"FFAD",x"FFAB",x"FFA5",x"FFA6",x"FFA7",x"FFAA",x"FFAA",x"FFB2",x"FFB7",x"FFC1",x"FFC9",x"FFD6",x"FFE0",x"FFEB",x"FFF8",x"0005",
    x"0014",x"0020",x"002C",x"0036",x"0043",x"004A",x"0053",x"005B",x"0061",x"0065",x"0068",x"006B",x"006C",x"006C",x"0068",x"0062",
    x"005F",x"0055",x"0050",x"0048",x"0042",x"0038",x"002E",x"0020",x"0018",x"000A",x"0005",x"FFF8",x"FFF0",x"FFE8",x"FFDD",x"FFD6",
    x"FFCF",x"FFCB",x"FFC8",x"FFC5",x"FFC3",x"FFC6",x"FFC8",x"FFCD",x"FFD2",x"FFD8",x"FFDF",x"FFE5",x"FFEE",x"FFF5",x"FFFF",x"0008",
    x"000E",x"0016",x"001D",x"0026",x"002D",x"0032",x"0037",x"003C",x"0040",x"0040",x"0044",x"0042",x"0043",x"0040",x"003B",x"0037",
    x"0031",x"002D",x"0023",x"001E",x"0015",x"000B",x"FFFF",x"FFF7",x"FFEC",x"FFE4",x"FFDC",x"FFD4",x"FFCD",x"FFC7",x"FFC0",x"FFBA",
    x"FFB5",x"FFB4",x"FFB2",x"FFB0",x"FFAF",x"FFB2",x"FFB6",x"FFB7",x"FFBC",x"FFC2",x"FFC7",x"FFCE",x"FFD7",x"FFDD",x"FFE5",x"FFF0",
    x"FFF8",x"0002",x"000B",x"0014",x"001B",x"0023",x"002C",x"0031",x"0039",x"003C",x"0040",x"0043",x"0046",x"0046",x"0048",x"0046",
    x"0044",x"0041",x"003D",x"0035",x"0031",x"0029",x"0021",x"001B",x"0014",x"0009",x"0003",x"FFF7",x"FFF0",x"FFE9",x"FFE1",x"FFDB",
    x"FFD4",x"FFD0",x"FFCA",x"FFC6",x"FFC3",x"FFC1",x"FFC0",x"FFBE",x"FFBD",x"FFC0",x"FFC2",x"FFC7",x"FFCB",x"FFCF",x"FFD3",x"FFDA",
    x"FFDF",x"FFE6",x"FFED",x"FFF2",x"FFF9",x"0000",x"0004",x"000A",x"0011",x"0014",x"0019",x"001E",x"0020",x"0022",x"0024",x"0024",
    x"0027",x"0027",x"0025",x"0026",x"0024",x"0021",x"001D",x"001C",x"0019",x"0015",x"0012",x"000E",x"000A",x"0005",x"0002",x"FFFE",
    x"FFF8",x"FFF5",x"FFF3",x"FFEF",x"FFEC",x"FFEA",x"FFE9",x"FFE7",x"FFE6",x"FFE6",x"FFE7",x"FFE8",x"FFE9",x"FFEB",x"FFEB",x"FFED",
    x"FFF0",x"FFF1",x"FFF4",x"FFF6",x"FFF8",x"FFFB",x"FFFE",x"0002",x"0004",x"0006",x"0008",x"0009",x"000B",x"000A",x"000A",x"000A",
    x"000B",x"000B",x"000A",x"0008",x"0007",x"0005",x"0003",x"0000",x"0000",x"FFFD",x"FFFC",x"FFF9",x"FFF7",x"FFF6",x"FFF3",x"FFF2",
    x"FFEF",x"FFEE",x"FFEC",x"FFEB",x"FFE9",x"FFE8",x"FFE9",x"FFE8",x"FFEA",x"FFEA",x"FFEA",x"FFEC",x"FFEC",x"FFEF",x"FFF1",x"FFF2",
    x"FFF4",x"FFF6",x"FFF7",x"FFF9",x"FFFA",x"FFFD",x"FFFE",x"FFFF",x"0001",x"0002",x"0004",x"0003",x"0004",x"0005",x"0007",x"0007",
    x"0007",x"0008",x"0008",x"0008",x"0007",x"0006",x"0006",x"0006",x"0004",x"0003",x"0003",x"0002",x"0001",x"FFFF",x"FFFE",x"FFFE",
    x"FFFD",x"FFFC",x"FFFC",x"FFFC",x"FFFB",x"FFFB",x"FFFB",x"FFFC",x"FFFD",x"FFFD",x"FFFF",x"0000",x"0001",x"0002",x"0002",x"0003",
    x"0004",x"0004",x"0005",x"0006",x"0008",x"0008",x"0009",x"0009",x"000B",x"000B",x"000C",x"000C",x"000C",x"000B",x"000A",x"000A",
    x"0008",x"0007",x"0006",x"0003",x"0002",x"0000",x"FFFE",x"FFFD",x"FFFA",x"FFF9",x"FFF7",x"FFF6",x"FFF5",x"FFF4",x"FFF2",x"FFF1",
    x"FFF1",x"FFF1",x"FFF0",x"FFEF",x"FFEF",x"FFF0",x"FFEF",x"FFF0",x"FFF1",x"FFF2",x"FFF4",x"FFF5",x"FFF7",x"FFF8",x"FFFA",x"FFFC",
    x"FFFD",x"FFFE",x"0000",x"0002",x"0003",x"0004",x"0006",x"0006",x"0008",x"0008",x"000A",x"000B",x"000C",x"000C",x"000D",x"000D",
    x"000D",x"000D",x"000C",x"000C",x"000B",x"000B",x"000A",x"0009",x"0008",x"0006",x"0006",x"0004",x"0002",x"0001",x"0001",x"0000",
    x"FFFF",x"FFFE",x"FFFE",x"FFFD",x"FFFD",x"FFFD",x"FFFC",x"FFFC",x"FFFC",x"FFFC",x"FFFC",x"FFFC",x"FFFD",x"FFFD",x"FFFE",x"FFFE",
    x"FFFE",x"FFFE",x"FFFF",x"0000",x"0001",x"0001",x"0002",x"0002",x"0002",x"0003",x"0004",x"0004",x"0004",x"0004",x"0005",x"0005",
    x"0004",x"0004",x"0004",x"0003",x"0003",x"0002",x"0002",x"0002",x"0002",x"0001",x"0001",x"0001",x"0000",x"FFFF",x"FFFF",x"FFFE",
    x"FFFE",x"FFFE",x"FFFD",x"FFFD",x"FFFC",x"FFFC",x"FFFD",x"FFFD",x"FFFD",x"FFFD",x"FFFD",x"FFFD",x"FFFE",x"FFFE",x"FFFF",x"0000",
    x"0000",x"0001",x"0001",x"0001",x"0002",x"0002",x"0003",x"0003",x"0003",x"0003",x"0003",x"0003",x"0003",x"0003",x"0003",x"0003",
    x"0002",x"0002",x"0002",x"0002",x"0001",x"0000",x"0000",x"0000",x"FFFF",x"FFFE",x"FFFE",x"FFFD",x"FFFC",x"FFFC",x"FFFB",x"FFFA",
    x"FFFA",x"FFFA",x"FFFA",x"FFFA",x"FFF9",x"FFF9",x"FFF9",x"FFF9",x"FFF9",x"FFFA",x"FFFA",x"FFFA",x"FFFA",x"FFFB",x"FFFC",x"FFFD",
    x"FFFD",x"FFFE",x"FFFF",x"FFFF",x"0000",x"0001",x"0002",x"0002",x"0004",x"0004",x"0005",x"0005",x"0006",x"0006",x"0007",x"0007",
    x"0007",x"0008",x"0008",x"0008",x"0007",x"0007",x"0007",x"0007",x"0006",x"0006",x"0005",x"0005",x"0004",x"0003",x"0003",x"0002",
    x"0001",x"0001",x"0000",x"FFFF",x"FFFE",x"FFFE",x"FFFD",x"FFFC",x"FFFC",x"FFFB",x"FFFA",x"FFFA",x"FFF9",x"FFF9",x"FFF9",x"FFF9",
    x"FFF9",x"FFF9",x"FFF9",x"FFF9",x"FFFA",x"FFFA",x"FFFB",x"FFFB",x"FFFB",x"FFFC",x"FFFC",x"FFFD",x"FFFD",x"FFFE",x"FFFF",x"0000"
  );
begin
  process(clock) is
  begin
    if rising_edge(clock) then
      data0_1 <= sound_data(to_integer(unsigned(addr0_0)));
      data1_1 <= sound_data(to_integer(unsigned(addr1_0)));
    end if;
  end process;
end v1;
