----------------------------------------------------------------------------------------------------------------------------------------------------------------
-- LSD.TOS, March 2017 (DO NOT REMOVE THIS LINE)
--
-- 8x8 font (in bold face) with 128 characters.
--
-- Source (public domain):
--   Daniel Hepper and Marcel Sondaar
--   https://github.com/dhepper/font8x8
--   font8x8_basic.h
--
-- Modified, expanded to 128 characters, and converted to VHDL.
--

library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

entity font_8x8_bold is
  port
  (
    clock : in std_logic; -- main clock

    char_0   : in  std_logic_vector(6 downto 0); -- character number encoded as a std_logic_vector
    row_0    : in  std_logic_vector(2 downto 0); -- row number encoded as a std_logic_vector: 0 (top) to 7 (bottom)
    column_0 : in  std_logic_vector(2 downto 0); -- column number encoded as a std_logic_vector: 0 (left) to 7 (right)
    data_1   : out std_logic                     -- pixel color ('0' means background color, '1' means foreground color)
  );
end font_8x8_bold;

architecture v1 of font_8x8_bold is
  signal addr_0x : std_logic_vector(12 downto 0); -- equal to 64*char+8*row+col
  --
  -- Single port ROM memory data
  --
  type rom_t is array(0 to 128*8*8-1) of std_logic;
  constant font_data : rom_t :=
  -- [  0,"0000000",0x00] top-left of a table box
    "00000000" &
    "00000000" &
    "00000000" &
    "00011111" &
    "00011111" &
    "00011000" &
    "00011000" &
    "00011000" &
  -- [  1,"0000001",0x01] top-center of a table box
    "00000000" &
    "00000000" &
    "00000000" &
    "11111111" &
    "11111111" &
    "00011000" &
    "00011000" &
    "00011000" &
  -- [  2,"0000010",0x02] top-right of a table box
    "00000000" &
    "00000000" &
    "00000000" &
    "11111000" &
    "11111000" &
    "00011000" &
    "00011000" &
    "00011000" &
  -- [  3,"0000011",0x03] middle-left of a table box
    "00011000" &
    "00011000" &
    "00011000" &
    "00011111" &
    "00011111" &
    "00011000" &
    "00011000" &
    "00011000" &
  -- [  4,"0000100",0x04] middle-center of a table box
    "00011000" &
    "00011000" &
    "00011000" &
    "11111111" &
    "11111111" &
    "00011000" &
    "00011000" &
    "00011000" &
  -- [  5,"0000101",0x05] middle-right of a table box
    "00011000" &
    "00011000" &
    "00011000" &
    "11111000" &
    "11111000" &
    "00011000" &
    "00011000" &
    "00011000" &
  -- [  6,"0000110",0x06] bottom-left of a table box
    "00011000" &
    "00011000" &
    "00011000" &
    "00011111" &
    "00011111" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [  7,"0000111",0x07] bottom-center of a table box
    "00011000" &
    "00011000" &
    "00011000" &
    "11111111" &
    "11111111" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [  8,"0001000",0x08] bottom-right of a table box
    "00011000" &
    "00011000" &
    "00011000" &
    "11111000" &
    "11111000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [  9,"0001001",0x09] horizontal line of a table box
    "00000000" &
    "00000000" &
    "00000000" &
    "11111111" &
    "11111111" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 10,"0001010",0x0A] vertical line of a table box
    "00011000" &
    "00011000" &
    "00011000" &
    "00011000" &
    "00011000" &
    "00011000" &
    "00011000" &
    "00011000" &
  -- [ 11,"0001011",0x0B] rounded top-left of a table box
    "00000000" &
    "00000000" &
    "00000000" &
    "00001111" &
    "00011111" &
    "00011000" &
    "00011000" &
    "00011000" &
  -- [ 12,"0001100",0x0C] rounded top-right of a table box
    "00000000" &
    "00000000" &
    "00000000" &
    "11110000" &
    "11111000" &
    "00011000" &
    "00011000" &
    "00011000" &
  -- [ 13,"0001101",0x0D] rounded bottom-left of a table box
    "00011000" &
    "00011000" &
    "00011000" &
    "00011111" &
    "00001111" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 14,"0001110",0x0E] rounded bottom-right of a table box
    "00011000" &
    "00011000" &
    "00011000" &
    "11111000" &
    "11110000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 15,"0001111",0x0F] thin X inside a box
    "11111111" &
    "11000011" &
    "10100101" &
    "10011001" &
    "10011001" &
    "10100101" &
    "11000011" &
    "11111111" &
  -- [ 16,"0010000",0x10] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 17,"0010001",0x11] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 18,"0010010",0x12] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 19,"0010011",0x13] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 20,"0010100",0x14] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 21,"0010101",0x15] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 22,"0010110",0x16] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 23,"0010111",0x17] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 24,"0011000",0x18] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 25,"0011001",0x19] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 26,"0011010",0x1A] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 27,"0011011",0x1B] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 28,"0011100",0x1C] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 29,"0011101",0x1D] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 30,"0011110",0x1E] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 31,"0011111",0x1F] unused (blank)
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 32,"0100000",0x20] space
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 33,"0100001",0x21] !
    "00011000" &
    "00111100" &
    "00111100" &
    "00011000" &
    "00011000" &
    "00000000" &
    "00011000" &
    "00000000" &
  -- [ 34,"0100010",0x22] "
    "01101100" &
    "01101100" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 35,"0100011",0x23] #
    "01101100" &
    "01101100" &
    "11111110" &
    "01101100" &
    "11111110" &
    "01101100" &
    "01101100" &
    "00000000" &
  -- [ 36,"0100100",0x24] $
    "00110000" &
    "01111100" &
    "11000000" &
    "01111000" &
    "00001100" &
    "11111000" &
    "00110000" &
    "00000000" &
  -- [ 37,"0100101",0x25] %
    "00000000" &
    "11000110" &
    "11001100" &
    "00011000" &
    "00110000" &
    "01100110" &
    "11000110" &
    "00000000" &
  -- [ 38,"0100110",0x26] &
    "00111000" &
    "01101100" &
    "00111000" &
    "01110110" &
    "11011100" &
    "11001100" &
    "01110110" &
    "00000000" &
  -- [ 39,"0100111",0x27] '
    "00011000" &
    "00011000" &
    "00110000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 40,"0101000",0x28] (
    "00011000" &
    "00110000" &
    "01100000" &
    "01100000" &
    "01100000" &
    "00110000" &
    "00011000" &
    "00000000" &
  -- [ 41,"0101001",0x29] )
    "01100000" &
    "00110000" &
    "00011000" &
    "00011000" &
    "00011000" &
    "00110000" &
    "01100000" &
    "00000000" &
  -- [ 42,"0101010",0x2A] *
    "00000000" &
    "01100110" &
    "00111100" &
    "11111111" &
    "00111100" &
    "01100110" &
    "00000000" &
    "00000000" &
  -- [ 43,"0101011",0x2B] +
    "00000000" &
    "00110000" &
    "00110000" &
    "11111100" &
    "00110000" &
    "00110000" &
    "00000000" &
    "00000000" &
  -- [ 44,"0101100",0x2C] ,
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00110000" &
    "00110000" &
    "01100000" &
  -- [ 45,"0101101",0x2D] -
    "00000000" &
    "00000000" &
    "00000000" &
    "11111100" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 46,"0101110",0x2E] .
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00110000" &
    "00110000" &
    "00000000" &
  -- [ 47,"0101111",0x2F] /
    "00000110" &
    "00001100" &
    "00011000" &
    "00110000" &
    "01100000" &
    "11000000" &
    "10000000" &
    "00000000" &
  -- [ 48,"0110000",0x30] 0
    "01111100" &
    "11000110" &
    "11001110" &
    "11011110" &
    "11110110" &
    "11100110" &
    "01111100" &
    "00000000" &
  -- [ 49,"0110001",0x31] 1
    "00110000" &
    "01110000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "11111100" &
    "00000000" &
  -- [ 50,"0110010",0x32] 2
    "01111000" &
    "11001100" &
    "00001100" &
    "00111000" &
    "01100000" &
    "11001100" &
    "11111100" &
    "00000000" &
  -- [ 51,"0110011",0x33] 3
    "01111000" &
    "11001100" &
    "00001100" &
    "00111000" &
    "00001100" &
    "11001100" &
    "01111000" &
    "00000000" &
  -- [ 52,"0110100",0x34] 4
    "00011100" &
    "00111100" &
    "01101100" &
    "11001100" &
    "11111110" &
    "00001100" &
    "00011110" &
    "00000000" &
  -- [ 53,"0110101",0x35] 5
    "11111100" &
    "11000000" &
    "11111000" &
    "00001100" &
    "00001100" &
    "11001100" &
    "01111000" &
    "00000000" &
  -- [ 54,"0110110",0x36] 6
    "00111000" &
    "01100000" &
    "11000000" &
    "11111000" &
    "11001100" &
    "11001100" &
    "01111000" &
    "00000000" &
  -- [ 55,"0110111",0x37] 7
    "11111100" &
    "11001100" &
    "00001100" &
    "00011000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "00000000" &
  -- [ 56,"0111000",0x38] 8
    "01111000" &
    "11001100" &
    "11001100" &
    "01111000" &
    "11001100" &
    "11001100" &
    "01111000" &
    "00000000" &
  -- [ 57,"0111001",0x39] 9
    "01111000" &
    "11001100" &
    "11001100" &
    "01111100" &
    "00001100" &
    "00011000" &
    "01110000" &
    "00000000" &
  -- [ 58,"0111010",0x3A] :
    "00000000" &
    "00110000" &
    "00110000" &
    "00000000" &
    "00000000" &
    "00110000" &
    "00110000" &
    "00000000" &
  -- [ 59,"0111011",0x3B] ;
    "00000000" &
    "00110000" &
    "00110000" &
    "00000000" &
    "00000000" &
    "00110000" &
    "00110000" &
    "01100000" &
  -- [ 60,"0111100",0x3C] <
    "00011000" &
    "00110000" &
    "01100000" &
    "11000000" &
    "01100000" &
    "00110000" &
    "00011000" &
    "00000000" &
  -- [ 61,"0111101",0x3D] =
    "00000000" &
    "00000000" &
    "11111100" &
    "00000000" &
    "00000000" &
    "11111100" &
    "00000000" &
    "00000000" &
  -- [ 62,"0111110",0x3E] >
    "01100000" &
    "00110000" &
    "00011000" &
    "00001100" &
    "00011000" &
    "00110000" &
    "01100000" &
    "00000000" &
  -- [ 63,"0111111",0x3F] ?
    "01111000" &
    "11001100" &
    "00001100" &
    "00011000" &
    "00110000" &
    "00000000" &
    "00110000" &
    "00000000" &
  -- [ 64,"1000000",0x40] @
    "01111100" &
    "11000110" &
    "11011110" &
    "11011110" &
    "11011110" &
    "11000000" &
    "01111000" &
    "00000000" &
  -- [ 65,"1000001",0x41] A
    "00110000" &
    "01111000" &
    "11001100" &
    "11001100" &
    "11111100" &
    "11001100" &
    "11001100" &
    "00000000" &
  -- [ 66,"1000010",0x42] B
    "11111100" &
    "01100110" &
    "01100110" &
    "01111100" &
    "01100110" &
    "01100110" &
    "11111100" &
    "00000000" &
  -- [ 67,"1000011",0x43] C
    "00111100" &
    "01100110" &
    "11000000" &
    "11000000" &
    "11000000" &
    "01100110" &
    "00111100" &
    "00000000" &
  -- [ 68,"1000100",0x44] D
    "11111000" &
    "01101100" &
    "01100110" &
    "01100110" &
    "01100110" &
    "01101100" &
    "11111000" &
    "00000000" &
  -- [ 69,"1000101",0x45] E
    "11111110" &
    "01100010" &
    "01101000" &
    "01111000" &
    "01101000" &
    "01100010" &
    "11111110" &
    "00000000" &
  -- [ 70,"1000110",0x46] F
    "11111110" &
    "01100010" &
    "01101000" &
    "01111000" &
    "01101000" &
    "01100000" &
    "11110000" &
    "00000000" &
  -- [ 71,"1000111",0x47] G
    "00111100" &
    "01100110" &
    "11000000" &
    "11000000" &
    "11001110" &
    "01100110" &
    "00111110" &
    "00000000" &
  -- [ 72,"1001000",0x48] H
    "11001100" &
    "11001100" &
    "11001100" &
    "11111100" &
    "11001100" &
    "11001100" &
    "11001100" &
    "00000000" &
  -- [ 73,"1001001",0x49] I
    "01111000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "01111000" &
    "00000000" &
  -- [ 74,"1001010",0x4A] J
    "00011110" &
    "00001100" &
    "00001100" &
    "00001100" &
    "11001100" &
    "11001100" &
    "01111000" &
    "00000000" &
  -- [ 75,"1001011",0x4B] K
    "11100110" &
    "01100110" &
    "01101100" &
    "01111000" &
    "01101100" &
    "01100110" &
    "11100110" &
    "00000000" &
  -- [ 76,"1001100",0x4C] L
    "11110000" &
    "01100000" &
    "01100000" &
    "01100000" &
    "01100010" &
    "01100110" &
    "11111110" &
    "00000000" &
  -- [ 77,"1001101",0x4D] M
    "11000110" &
    "11101110" &
    "11111110" &
    "11111110" &
    "11010110" &
    "11000110" &
    "11000110" &
    "00000000" &
  -- [ 78,"1001110",0x4E] N
    "11000110" &
    "11100110" &
    "11110110" &
    "11011110" &
    "11001110" &
    "11000110" &
    "11000110" &
    "00000000" &
  -- [ 79,"1001111",0x4F] O
    "00111000" &
    "01101100" &
    "11000110" &
    "11000110" &
    "11000110" &
    "01101100" &
    "00111000" &
    "00000000" &
  -- [ 80,"1010000",0x50] P
    "11111100" &
    "01100110" &
    "01100110" &
    "01111100" &
    "01100000" &
    "01100000" &
    "11110000" &
    "00000000" &
  -- [ 81,"1010001",0x51] Q
    "01111000" &
    "11001100" &
    "11001100" &
    "11001100" &
    "11011100" &
    "01111000" &
    "00011100" &
    "00000000" &
  -- [ 82,"1010010",0x52] R
    "11111100" &
    "01100110" &
    "01100110" &
    "01111100" &
    "01101100" &
    "01100110" &
    "11100110" &
    "00000000" &
  -- [ 83,"1010011",0x53] S
    "01111000" &
    "11001100" &
    "11100000" &
    "01110000" &
    "00011100" &
    "11001100" &
    "01111000" &
    "00000000" &
  -- [ 84,"1010100",0x54] T
    "11111100" &
    "10110100" &
    "00110000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "01111000" &
    "00000000" &
  -- [ 85,"1010101",0x55] U
    "11001100" &
    "11001100" &
    "11001100" &
    "11001100" &
    "11001100" &
    "11001100" &
    "11111100" &
    "00000000" &
  -- [ 86,"1010110",0x56] V
    "11001100" &
    "11001100" &
    "11001100" &
    "11001100" &
    "11001100" &
    "01111000" &
    "00110000" &
    "00000000" &
  -- [ 87,"1010111",0x57] W
    "11000110" &
    "11000110" &
    "11000110" &
    "11010110" &
    "11111110" &
    "11101110" &
    "11000110" &
    "00000000" &
  -- [ 88,"1011000",0x58] X
    "11000110" &
    "11000110" &
    "01101100" &
    "00111000" &
    "00111000" &
    "01101100" &
    "11000110" &
    "00000000" &
  -- [ 89,"1011001",0x59] Y
    "11001100" &
    "11001100" &
    "11001100" &
    "01111000" &
    "00110000" &
    "00110000" &
    "01111000" &
    "00000000" &
  -- [ 90,"1011010",0x5A] Z
    "11111110" &
    "11000110" &
    "10001100" &
    "00011000" &
    "00110010" &
    "01100110" &
    "11111110" &
    "00000000" &
  -- [ 91,"1011011",0x5B] [
    "01111000" &
    "01100000" &
    "01100000" &
    "01100000" &
    "01100000" &
    "01100000" &
    "01111000" &
    "00000000" &
  -- [ 92,"1011100",0x5C] \
    "11000000" &
    "01100000" &
    "00110000" &
    "00011000" &
    "00001100" &
    "00000110" &
    "00000010" &
    "00000000" &
  -- [ 93,"1011101",0x5D] ]
    "01111000" &
    "00011000" &
    "00011000" &
    "00011000" &
    "00011000" &
    "00011000" &
    "01111000" &
    "00000000" &
  -- [ 94,"1011110",0x5E] ^
    "00010000" &
    "00111000" &
    "01101100" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 95,"1011111",0x5F] _
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "11111110" &
  -- [ 96,"1100000",0x60] `
    "00110000" &
    "00110000" &
    "00011000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [ 97,"1100001",0x61] a
    "00000000" &
    "00000000" &
    "01111000" &
    "00001100" &
    "01111100" &
    "11001100" &
    "01110110" &
    "00000000" &
  -- [ 98,"1100010",0x62] b
    "11100000" &
    "01100000" &
    "01100000" &
    "01111100" &
    "01100110" &
    "01100110" &
    "11011100" &
    "00000000" &
  -- [ 99,"1100011",0x63] c
    "00000000" &
    "00000000" &
    "01111000" &
    "11001100" &
    "11000000" &
    "11001100" &
    "01111000" &
    "00000000" &
  -- [100,"1100100",0x64] d
    "00011100" &
    "00001100" &
    "00001100" &
    "01111100" &
    "11001100" &
    "11001100" &
    "01110110" &
    "00000000" &
  -- [101,"1100101",0x65] e
    "00000000" &
    "00000000" &
    "01111000" &
    "11001100" &
    "11111100" &
    "11000000" &
    "01111000" &
    "00000000" &
  -- [102,"1100110",0x66] f
    "00111000" &
    "01101100" &
    "01100000" &
    "11110000" &
    "01100000" &
    "01100000" &
    "11110000" &
    "00000000" &
  -- [103,"1100111",0x67] g
    "00000000" &
    "00000000" &
    "01110110" &
    "11001100" &
    "11001100" &
    "01111100" &
    "00001100" &
    "11111000" &
  -- [104,"1101000",0x68] h
    "11100000" &
    "01100000" &
    "01101100" &
    "01110110" &
    "01100110" &
    "01100110" &
    "11100110" &
    "00000000" &
  -- [105,"1101001",0x69] i
    "00110000" &
    "00000000" &
    "01110000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "01111000" &
    "00000000" &
  -- [106,"1101010",0x6A] j
    "00001100" &
    "00000000" &
    "00001100" &
    "00001100" &
    "00001100" &
    "11001100" &
    "11001100" &
    "01111000" &
  -- [107,"1101011",0x6B] k
    "11100000" &
    "01100000" &
    "01100110" &
    "01101100" &
    "01111000" &
    "01101100" &
    "11100110" &
    "00000000" &
  -- [108,"1101100",0x6C] l
    "01110000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "00110000" &
    "01111000" &
    "00000000" &
  -- [109,"1101101",0x6D] m
    "00000000" &
    "00000000" &
    "11001100" &
    "11111110" &
    "11111110" &
    "11010110" &
    "11000110" &
    "00000000" &
  -- [110,"1101110",0x6E] n
    "00000000" &
    "00000000" &
    "11111000" &
    "11001100" &
    "11001100" &
    "11001100" &
    "11001100" &
    "00000000" &
  -- [111,"1101111",0x6F] o
    "00000000" &
    "00000000" &
    "01111000" &
    "11001100" &
    "11001100" &
    "11001100" &
    "01111000" &
    "00000000" &
  -- [112,"1110000",0x70] p
    "00000000" &
    "00000000" &
    "11011100" &
    "01100110" &
    "01100110" &
    "01111100" &
    "01100000" &
    "11110000" &
  -- [113,"1110001",0x71] q
    "00000000" &
    "00000000" &
    "01110110" &
    "11001100" &
    "11001100" &
    "01111100" &
    "00001100" &
    "00011110" &
  -- [114,"1110010",0x72] r
    "00000000" &
    "00000000" &
    "11011100" &
    "01110110" &
    "01100110" &
    "01100000" &
    "11110000" &
    "00000000" &
  -- [115,"1110011",0x73] s
    "00000000" &
    "00000000" &
    "01111100" &
    "11000000" &
    "01111000" &
    "00001100" &
    "11111000" &
    "00000000" &
  -- [116,"1110100",0x74] t
    "00010000" &
    "00110000" &
    "01111100" &
    "00110000" &
    "00110000" &
    "00110100" &
    "00011000" &
    "00000000" &
  -- [117,"1110101",0x75] u
    "00000000" &
    "00000000" &
    "11001100" &
    "11001100" &
    "11001100" &
    "11001100" &
    "01110110" &
    "00000000" &
  -- [118,"1110110",0x76] v
    "00000000" &
    "00000000" &
    "11001100" &
    "11001100" &
    "11001100" &
    "01111000" &
    "00110000" &
    "00000000" &
  -- [119,"1110111",0x77] w
    "00000000" &
    "00000000" &
    "11000110" &
    "11010110" &
    "11111110" &
    "11111110" &
    "01101100" &
    "00000000" &
  -- [120,"1111000",0x78] x
    "00000000" &
    "00000000" &
    "11000110" &
    "01101100" &
    "00111000" &
    "01101100" &
    "11000110" &
    "00000000" &
  -- [121,"1111001",0x79] y
    "00000000" &
    "00000000" &
    "11001100" &
    "11001100" &
    "11001100" &
    "01111100" &
    "00001100" &
    "11111000" &
  -- [122,"1111010",0x7A] z
    "00000000" &
    "00000000" &
    "11111100" &
    "10011000" &
    "00110000" &
    "01100100" &
    "11111100" &
    "00000000" &
  -- [123,"1111011",0x7B] {
    "00011100" &
    "00110000" &
    "00110000" &
    "11100000" &
    "00110000" &
    "00110000" &
    "00011100" &
    "00000000" &
  -- [124,"1111100",0x7C] |
    "00011000" &
    "00011000" &
    "00011000" &
    "00000000" &
    "00011000" &
    "00011000" &
    "00011000" &
    "00000000" &
  -- [125,"1111101",0x7D] }
    "11100000" &
    "00110000" &
    "00110000" &
    "00011100" &
    "00110000" &
    "00110000" &
    "11100000" &
    "00000000" &
  -- [126,"1111110",0x7E] ~
    "01110110" &
    "11011100" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
    "00000000" &
  -- [127,"1111111",0x7F] filled o (a disk)
    "00000000" &
    "00000000" &
    "01111000" &
    "11111100" &
    "11111100" &
    "11111100" &
    "01111000" &
    "00000000";
begin
  addr_0x <= char_0 & row_0 & column_0;
  process(clock) is
  begin
    if rising_edge(clock) then
      data_1 <= font_data(to_integer(unsigned(addr_0x)));
    end if;
  end process;
end v1;
