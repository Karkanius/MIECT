library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity ROM_sin is
	port(address	: in  std_logic_vector(7 downto 0);
		  sin_out	: out std_logic_vector(15 downto 0));
end ROM_sin;

architecture Behavioral of ROM_sin is
	
	type sin is array (0 to 255) of integer;
	constant sin1 : sin := (0, 807, 1614, 2419, 3224, 4026, 4826, 5623, 6417, 7207, 7992, 8772,
									9548, 10317, 11080, 11836, 12586, 13327, 14061, 14786, 15502, 16208,
									16905, 17591, 18267, 18932, 19585, 20226, 20855, 21472, 22075, 22665,
									23241, 23803, 24350, 24883, 25401, 25903, 26390, 26860, 27315, 27752,
									28173, 28577, 28963, 29332, 29683, 30016, 30330, 30627, 30904, 31163,
									31403, 31624, 31826, 32008, 32171, 32315, 32439, 32543, 32627, 32692,
									32737, 32761, 32766, 32751, 32717, 32662, 32587, 32493, 32379, 32246,
									32092, 31920, 31727, 31516, 31286, 31036, 30768, 30481, 30175, 29851,
									29509, 29150, 28772, 28377, 27965, 27535, 27090, 26627, 26149, 25654,
									25144, 24619, 24079, 23524, 22955, 22371, 21775, 21165, 20542, 19907,
									19260, 18601, 17931, 17249, 16558, 15856, 15145, 14424, 13695, 12957,
									12212, 11459, 10699, 9933, 9161, 8383, 7600, 6812, 6021, 5225, 4427,
									3625, 2822, 2017, 1210, 403, -403, -1210, -2017, -2822, -3625, -4427,
									-5225, -6021, -6812, -7600, -8383, -9161, -9933, -10699, -11459, -12212,
									-12957, -13695, -14424, -15145, -15856, -16558, -17249, -17931, -18601,
									-19260, -19907, -20542, -21165, -21775, -22371, -22955, -23524, -24079,
									-24619, -25144, -25654, -26149, -26627, -27090, -27535, -27965, -28377,
									-28772, -29150, -29509, -29851, -30175, -30481, -30768, -31036, -31286,
									-31516, -31727, -31920, -32092, -32246, -32379, -32493, -32587, -32662,
									-32717, -32751, -32766, -32761, -32737, -32692, -32627, -32543, -32439,
									-32315, -32171, -32008, -31826, -31624, -31403, -31163, -30904, -30627,
									-30330, -30016, -29683, -29332, -28963, -28577, -28173, -27752, -27315,
									-26860, -26390, -25903, -25401, -24883, -24350, -23803, -23241, -22665,
									-22075, -21472, -20855, -20226, -19585, -18932, -18267, -17591, -16905,
									-16208, -15502, -14786, -14061, -13327, -12586, -11836, -11080, -10317,
									-9548, -8772, -7992, -7207, -6417, -5623, -4826, -4026, -3224, -2419,
									-1614, -807, 0);

begin
	sin_out <= std_logic_vector(to_signed(sin1(to_integer(unsigned(address))), 16));
end Behavioral;
