--
--
--
--import java.util.*;
--
--public class FreqObtainer {
--	
--	public static void main (String[] args) {
--		
--		//Variáveis
--		double freq [] = { 261.63, 277.18, 293.66, 311.13, 329.63, 349.23, 369.99, 392.00, 415.30, 440.00, 466.16, 493.88, 0.00, 0.00, 0.00, 0.00 };
--		double fator;
--		
--		for (int i = 0; i < 16; i++)
--		{
--			System.out.printf("    -- nota %02d\n",i);
--			fator = 2.0 * Math.PI * freq[i] / 48000.0;
--			for(int j = 0; j < 1024; j++)
--			{
--				System.out.printf("    x\"%04X\",\n",0xFFFF & Math.round(32767.0 * Math.sin(fator*j)));
--			}
--		}
--		
--	}
--}
--
--
--
--
--
--Função escrita em java que permitiu o cálculo dos valores presentes nesta mesma ROM
--
--Mais detalhes no relatório enviado em anexo
--
--

library ieee;
use     ieee.std_logic_1164.all;
use     ieee.numeric_std.all;

entity sound_rom is
  port
  (
    clock   : in  std_logic;
    nota    : in  std_logic_vector( 3 downto 0);
    counter : in  std_logic_vector( 9 downto 0);
    sample  : out std_logic_vector(15 downto 0)
  );
end sound_rom;

architecture v1 of sound_rom is

  signal addr : std_logic_vector(13 downto 0);
  type rom_t is array(0 to 16*1024-1) of std_logic_vector(15 downto 0);
  
  constant rom : rom_t :=(
	    -- nota 00
    x"0000",
    x"08C3",
    x"117B",
    x"1A1E",
    x"22A2",
    x"2AFC",
    x"3322",
    x"3B0B",
    x"42AE",
    x"4A00",
    x"50F9",
    x"5792",
    x"5DC1",
    x"637F",
    x"68C6",
    x"6D8F",
    x"71D5",
    x"7592",
    x"78C2",
    x"7B61",
    x"7D6C",
    x"7EE0",
    x"7FBC",
    x"7FFF",
    x"7FA8",
    x"7EB7",
    x"7D2F",
    x"7B10",
    x"785D",
    x"751A",
    x"714B",
    x"6CF3",
    x"6819",
    x"62C1",
    x"5CF3",
    x"56B6",
    x"5010",
    x"490A",
    x"41AD",
    x"3A01",
    x"320F",
    x"29E1",
    x"2180",
    x"18F8",
    x"1051",
    x"0797",
    x"FED4",
    x"F612",
    x"ED5C",
    x"E4BD",
    x"DC3E",
    x"D3EA",
    x"CBCB",
    x"C3EB",
    x"BC53",
    x"B50C",
    x"AE1F",
    x"A794",
    x"A174",
    x"9BC5",
    x"968F",
    x"91D7",
    x"8DA3",
    x"89F8",
    x"86DC",
    x"8450",
    x"825A",
    x"80FA",
    x"8032",
    x"8004",
    x"8070",
    x"8175",
    x"8311",
    x"8544",
    x"880A",
    x"8B60",
    x"8F42",
    x"93AC",
    x"9897",
    x"9DFF",
    x"A3DC",
    x"AA28",
    x"B0DB",
    x"B7ED",
    x"BF55",
    x"C70B",
    x"CF06",
    x"D73B",
    x"DFA2",
    x"E82F",
    x"F0D9",
    x"F994",
    x"0258",
    x"0B19",
    x"13CC",
    x"1C68",
    x"24E2",
    x"2D2F",
    x"3546",
    x"3D1D",
    x"44AB",
    x"4BE6",
    x"52C7",
    x"5944",
    x"5F55",
    x"64F4",
    x"6A1A",
    x"6EC1",
    x"72E3",
    x"767A",
    x"7984",
    x"7BFC",
    x"7DDE",
    x"7F2A",
    x"7FDD",
    x"7FF6",
    x"7F76",
    x"7E5D",
    x"7CAC",
    x"7A66",
    x"778C",
    x"7423",
    x"702F",
    x"6BB4",
    x"66B7",
    x"613F",
    x"5B53",
    x"54F9",
    x"4E39",
    x"471A",
    x"3FA7",
    x"37E7",
    x"2FE4",
    x"27A8",
    x"1F3C",
    x"16AA",
    x"0DFD",
    x"0540",
    x"FC7C",
    x"F3BC",
    x"EB0B",
    x"E274",
    x"D9FF",
    x"D1B9",
    x"C9A9",
    x"C1DC",
    x"BA58",
    x"B329",
    x"AC55",
    x"A5E6",
    x"9FE4",
    x"9A54",
    x"953F",
    x"90AA",
    x"8C9A",
    x"8915",
    x"861F",
    x"83BB",
    x"81ED",
    x"80B5",
    x"8017",
    x"8012",
    x"80A6",
    x"81D4",
    x"8399",
    x"85F3",
    x"88E0",
    x"8C5C",
    x"9063",
    x"94F0",
    x"99FD",
    x"9F85",
    x"A580",
    x"ABE9",
    x"B2B6",
    x"B9E0",
    x"C15E",
    x"C927",
    x"D133",
    x"D976",
    x"E1E8",
    x"EA7D",
    x"F32D",
    x"FBEC",
    x"04B0",
    x"0D6E",
    x"161C",
    x"1EB0",
    x"271F",
    x"2F5F",
    x"3766",
    x"3F2A",
    x"46A3",
    x"4DC6",
    x"548D",
    x"5AEE",
    x"60E2",
    x"6661",
    x"6B66",
    x"6FE9",
    x"73E6",
    x"7758",
    x"7A3B",
    x"7C8B",
    x"7E46",
    x"7F69",
    x"7FF3",
    x"7FE3",
    x"7F3A",
    x"7DF8",
    x"7C1F",
    x"79B1",
    x"76B1",
    x"7322",
    x"6F09",
    x"6A6B",
    x"654D",
    x"5FB5",
    x"59AA",
    x"5334",
    x"4C5A",
    x"4524",
    x"3D9C",
    x"35C9",
    x"2DB6",
    x"256B",
    x"1CF4",
    x"145B",
    x"0BA8",
    x"02E8",
    x"FA24",
    x"F167",
    x"E8BC",
    x"E02D",
    x"D7C4",
    x"CF8B",
    x"C78C",
    x"BFD2",
    x"B864",
    x"B14C",
    x"AA93",
    x"A440",
    x"9E5B",
    x"98EC",
    x"93F8",
    x"8F86",
    x"8B9C",
    x"883C",
    x"856D",
    x"8331",
    x"818A",
    x"807C",
    x"8006",
    x"802B",
    x"80E8",
    x"823E",
    x"842C",
    x"86AD",
    x"89C1",
    x"8D62",
    x"918E",
    x"963D",
    x"9B6C",
    x"A113",
    x"A72D",
    x"ADB1",
    x"B498",
    x"BBD9",
    x"C36C",
    x"CB48",
    x"D363",
    x"DBB4",
    x"E430",
    x"ECCE",
    x"F583",
    x"FE44",
    x"0708",
    x"0FC3",
    x"186B",
    x"20F5",
    x"2959",
    x"318A",
    x"3980",
    x"4131",
    x"4894",
    x"4FA0",
    x"564C",
    x"5C90",
    x"6266",
    x"67C5",
    x"6CA7",
    x"7108",
    x"74E0",
    x"782C",
    x"7AE8",
    x"7D10",
    x"7EA3",
    x"7F9D",
    x"7FFE",
    x"7FC5",
    x"7EF3",
    x"7D88",
    x"7B87",
    x"78F2",
    x"75CB",
    x"7217",
    x"6DDA",
    x"6919",
    x"63D9",
    x"5E22",
    x"57FA",
    x"5169",
    x"4A75",
    x"4328",
    x"3B8B",
    x"33A6",
    x"2B83",
    x"232C",
    x"1AAB",
    x"1209",
    x"0952",
    x"0090",
    x"F7CD",
    x"EF14",
    x"E66F",
    x"DDE9",
    x"D58C",
    x"CD62",
    x"C574",
    x"BDCD",
    x"B676",
    x"AF76",
    x"A8D8",
    x"A2A2",
    x"9CDC",
    x"978D",
    x"92BB",
    x"8E6D",
    x"8AA7",
    x"876E",
    x"84C5",
    x"82B1",
    x"8133",
    x"804D",
    x"8001",
    x"804E",
    x"8135",
    x"82B4",
    x"84C9",
    x"8772",
    x"8AAC",
    x"8E73",
    x"92C2",
    x"9794",
    x"9CE3",
    x"A2AA",
    x"A8E1",
    x"AF80",
    x"B680",
    x"BDD8",
    x"C57F",
    x"CD6D",
    x"D598",
    x"DDF5",
    x"E67B",
    x"EF20",
    x"F7D9",
    x"009C",
    x"095E",
    x"1215",
    x"1AB7",
    x"2338",
    x"2B8F",
    x"33B1",
    x"3B96",
    x"4333",
    x"4A7F",
    x"5172",
    x"5803",
    x"5E2B",
    x"63E1",
    x"6920",
    x"6DE0",
    x"721C",
    x"75D0",
    x"78F6",
    x"7B8A",
    x"7D8B",
    x"7EF4",
    x"7FC6",
    x"7FFE",
    x"7F9C",
    x"7EA1",
    x"7D0E",
    x"7AE5",
    x"7828",
    x"74DB",
    x"7102",
    x"6CA1",
    x"67BE",
    x"625E",
    x"5C88",
    x"5643",
    x"4F96",
    x"488A",
    x"4127",
    x"3975",
    x"317F",
    x"294D",
    x"20E9",
    x"185E",
    x"0FB6",
    x"06FB",
    x"FE38",
    x"F576",
    x"ECC2",
    x"E424",
    x"DBA8",
    x"D358",
    x"CB3D",
    x"C361",
    x"BBCE",
    x"B48E",
    x"ADA7",
    x"A724",
    x"A10B",
    x"9B64",
    x"9636",
    x"9187",
    x"8D5D",
    x"89BC",
    x"86AA",
    x"8429",
    x"823C",
    x"80E7",
    x"802A",
    x"8007",
    x"807D",
    x"818C",
    x"8334",
    x"8571",
    x"8841",
    x"8BA1",
    x"8F8C",
    x"93FF",
    x"98F3",
    x"9E63",
    x"A449",
    x"AA9C",
    x"B156",
    x"B86E",
    x"BFDC",
    x"C798",
    x"CF97",
    x"D7D0",
    x"E039",
    x"E8C8",
    x"F174",
    x"FA31",
    x"02F4",
    x"0BB5",
    x"1467",
    x"1D00",
    x"2577",
    x"2DC1",
    x"35D4",
    x"3DA6",
    x"452F",
    x"4C64",
    x"533E",
    x"59B3",
    x"5FBD",
    x"6554",
    x"6A71",
    x"6F0F",
    x"7327",
    x"76B5",
    x"79B5",
    x"7C22",
    x"7DFA",
    x"7F3B",
    x"7FE4",
    x"7FF2",
    x"7F68",
    x"7E44",
    x"7C88",
    x"7A38",
    x"7754",
    x"73E1",
    x"6FE3",
    x"6B5F",
    x"665A",
    x"60D9",
    x"5AE5",
    x"5484",
    x"4DBD",
    x"4698",
    x"3F1F",
    x"375A",
    x"2F53",
    x"2713",
    x"1EA4",
    x"1610",
    x"0D62",
    x"04A4",
    x"FBE0",
    x"F321",
    x"EA71",
    x"E1DC",
    x"D96A",
    x"D127",
    x"C91C",
    x"C153",
    x"B9D5",
    x"B2AC",
    x"ABDF",
    x"A578",
    x"9F7D",
    x"99F6",
    x"94E9",
    x"905D",
    x"8C57",
    x"88DC",
    x"85F0",
    x"8396",
    x"81D2",
    x"80A5",
    x"8011",
    x"8017",
    x"80B7",
    x"81EF",
    x"83BE",
    x"8623",
    x"891A",
    x"8CA0",
    x"90B0",
    x"9546",
    x"9A5C",
    x"9FEC",
    x"A5EF",
    x"AC5F",
    x"B333",
    x"BA63",
    x"C1E6",
    x"C9B5",
    x"D1C4",
    x"DA0B",
    x"E280",
    x"EB18",
    x"F3C9",
    x"FC88",
    x"054C",
    x"0E0A",
    x"16B6",
    x"1F48",
    x"27B3",
    x"2FF0",
    x"37F2",
    x"3FB2",
    x"4725",
    x"4E42",
    x"5502",
    x"5B5B",
    x"6147",
    x"66BE",
    x"6BBA",
    x"7035",
    x"7428",
    x"7791",
    x"7A69",
    x"7CAF",
    x"7E5F",
    x"7F77",
    x"7FF7",
    x"7FDC",
    x"7F29",
    x"7DDC",
    x"7BF8",
    x"7980",
    x"7676",
    x"72DD",
    x"6EBB",
    x"6A14",
    x"64ED",
    x"5F4D",
    x"593B",
    x"52BD",
    x"4BDD",
    x"44A1",
    x"3D13",
    x"353B",
    x"2D24",
    x"24D6",
    x"1C5C",
    x"13C0",
    x"0B0D",
    x"024C",
    x"F988",
    x"F0CC",
    x"E823",
    x"DF96",
    x"D730",
    x"CEFB",
    x"C700",
    x"BF4B",
    x"B7E3",
    x"B0D1",
    x"AA1F",
    x"A3D3",
    x"9DF7",
    x"9890",
    x"93A5",
    x"8F3C",
    x"8B5B",
    x"8806",
    x"8540",
    x"830F",
    x"8173",
    x"806F",
    x"8004",
    x"8033",
    x"80FB",
    x"825C",
    x"8454",
    x"86E0",
    x"89FD",
    x"8DA8",
    x"91DD",
    x"9696",
    x"9BCD",
    x"A17C",
    x"A79D",
    x"AE29",
    x"B516",
    x"BC5D",
    x"C3F6",
    x"CBD6",
    x"D3F6",
    x"DC4A",
    x"E4C9",
    x"ED68",
    x"F61E",
    x"FEE0",
    x"07A3",
    x"105E",
    x"1904",
    x"218C",
    x"29EC",
    x"321A",
    x"3A0C",
    x"41B8",
    x"4915",
    x"501A",
    x"56BF",
    x"5CFC",
    x"62C9",
    x"6820",
    x"6CFA",
    x"7151",
    x"751F",
    x"7862",
    x"7B13",
    x"7D31",
    x"7EB9",
    x"7FA8",
    x"7FFF",
    x"7FBB",
    x"7EDF",
    x"7D69",
    x"7B5E",
    x"78BE",
    x"758D",
    x"71D0",
    x"6D89",
    x"68BF",
    x"6377",
    x"5DB8",
    x"5789",
    x"50F0",
    x"49F6",
    x"42A3",
    x"3B01",
    x"3317",
    x"2AF0",
    x"2296",
    x"1A12",
    x"116E",
    x"08B6",
    x"FFF4",
    x"F731",
    x"EE79",
    x"E5D6",
    x"DD53",
    x"D4F9",
    x"CCD2",
    x"C4EA",
    x"BD48",
    x"B5F6",
    x"AEFD",
    x"A865",
    x"A237",
    x"9C79",
    x"9733",
    x"926A",
    x"8E25",
    x"8A69",
    x"873A",
    x"849C",
    x"8292",
    x"811E",
    x"8043",
    x"8001",
    x"8059",
    x"814B",
    x"82D4",
    x"84F3",
    x"87A7",
    x"8AEB",
    x"8EBB",
    x"9313",
    x"97EE",
    x"9D47",
    x"A315",
    x"A953",
    x"AFF9",
    x"B700",
    x"BE5E",
    x"C60A",
    x"CDFD",
    x"D62B",
    x"DE8C",
    x"E714",
    x"EFBB",
    x"F875",
    x"0138",
    x"09FA",
    x"12B0",
    x"1B4F",
    x"23CE",
    x"2C22",
    x"3440",
    x"3C20",
    x"43B8",
    x"4AFE",
    x"51EA",
    x"5874",
    x"5E94",
    x"6443",
    x"6978",
    x"6E30",
    x"7263",
    x"760C",
    x"7928",
    x"7BB3",
    x"7DA9",
    x"7F08",
    x"7FCF",
    x"7FFC",
    x"7F8F",
    x"7E8A",
    x"7CEC",
    x"7AB9",
    x"77F2",
    x"749B",
    x"70B8",
    x"6C4E",
    x"6762",
    x"61F9",
    x"5C1C",
    x"55CF",
    x"4F1B",
    x"4809",
    x"40A0",
    x"38E9",
    x"30EF",
    x"28B9",
    x"2052",
    x"17C5",
    x"0F1B",
    x"065F",
    x"FD9C",
    x"F4DB",
    x"EC27",
    x"E38C",
    x"DB12",
    x"D2C5",
    x"CAAF",
    x"C2D8",
    x"BB4A",
    x"B410",
    x"AD30",
    x"A6B4",
    x"A0A3",
    x"9B04",
    x"95DF",
    x"9139",
    x"8D18",
    x"8981",
    x"8678",
    x"8401",
    x"821F",
    x"80D5",
    x"8023",
    x"800A",
    x"808B",
    x"81A5",
    x"8357",
    x"859E",
    x"8878",
    x"8BE2",
    x"8FD7",
    x"9453",
    x"9950",
    x"9EC9",
    x"A4B6",
    x"AB11",
    x"B1D1",
    x"B8F0",
    x"C064",
    x"C824",
    x"D027",
    x"D864",
    x"E0D0",
    x"E962",
    x"F20F",
    x"FACD",
    x"0390",
    x"0C50",
    x"1501",
    x"1D98",
    x"260D",
    x"2E53",
    x"3662",
    x"3E2F",
    x"45B2",
    x"4CE1",
    x"53B4",
    x"5A22",
    x"6025",
    x"65B3",
    x"6AC8",
    x"6F5C",
    x"736B",
    x"76EF",
    x"79E5",
    x"7C48",
    x"7E16",
    x"7F4C",
    x"7FEA",
    x"7FEE",
    x"7F58",
    x"7E2A",
    x"7C64",
    x"7A09",
    x"771B",
    x"739E",
    x"6F97",
    x"6B09",
    x"65FB",
    x"6073",
    x"5A77",
    x"540E",
    x"4D40",
    x"4616",
    x"3E97",
    x"36CD",
    x"2EC2",
    x"267E",
    x"1E0C",
    x"1576",
    x"0CC7",
    x"0408",
    x"FB44",
    x"F285",
    x"E9D7",
    x"E144",
    x"D8D5",
    x"D096",
    x"C88F",
    x"C0CB",
    x"B953",
    x"B230",
    x"AB6A",
    x"A50A",
    x"9F16",
    x"9998",
    x"9494",
    x"9011",
    x"8C14",
    x"88A3",
    x"85C1",
    x"8372",
    x"81B8",
    x"8096",
    x"800D",
    x"801D",
    x"80C7",
    x"820A",
    x"83E4",
    x"8653",
    x"8954",
    x"8CE4",
    x"90FD",
    x"959C",
    x"9ABB",
    x"A053",
    x"A65E",
    x"ACD5",
    x"B3B0",
    x"BAE6",
    x"C26F",
    x"CA42",
    x"D256",
    x"DAA0",
    x"E318",
    x"EBB2",
    x"F464",
    x"FD24",
    x"05E8",
    x"0EA5",
    x"1750",
    x"1FDF",
    x"2848",
    x"3080",
    x"387F",
    x"4039",
    x"47A6",
    x"4EBE",
    x"5576",
    x"5BC9",
    x"61AD",
    x"671B",
    x"6C0E",
    x"707F",
    x"746A",
    x"77C8",
    x"7A97",
    x"7CD2",
    x"7E77",
    x"7F85",
    x"7FFA",
    x"7FD5",
    x"7F16",
    x"7DBF",
    x"7BD1",
    x"794F",
    x"763A",
    x"7298",
    x"6E6C",
    x"69BC",
    x"648C",
    x"5EE4",
    x"58CA",
    x"5246",
    x"4B5F",
    x"441D",
    x"3C89",
    x"34AD",
    x"2C91",
    x"2440",
    x"1BC4",
    x"1326",
    x"0A71",
    x"01B0",
    x"F8EC",
    x"F031",
    x"E789",
    x"DEFF",
    x"D69C",
    x"CE6A",
    x"C675",
    x"BEC4",
    x"B762",
    x"B057",
    x"A9AB",
    x"A367",
    x"9D93",
    x"9834",
    x"9352",
    x"8EF3",
    x"8B1B",
    x"87D0",
    x"8514",
    x"82ED",
    x"815C",
    x"8062",
    x"8002",
    x"803C",
    x"810F",
    x"827A",
    x"847C",
    x"8712",
    x"8A3A",
    x"8DEF",
    x"922D",
    x"96EE",
    x"9C2E",
    x"A1E6",
    x"A80F",
    x"AEA1",
    x"B595",
    x"BCE2",
    x"C480",
    x"CC65",
    x"D488",
    x"DCE0",
    x"E562",
    x"EE03",
    x"F6BA",
    x"FF7C",
    x"083F",
    x"10F8",
    x"199D",
    x"2223",
    x"2A80",
    x"32AA",
    x"3A97",
    x"423D",
    x"4995",
    x"5093",
    x"5732",
    x"5D67",
    x"632C",
    x"687A",
    -- nota 01
    x"0000",
    x"0948",
    x"1283",
    x"1BA5",
    x"24A2",
    x"2D6E",
    x"35FC",
    x"3E42",
    x"4633",
    x"4DC7",
    x"54F1",
    x"5BA9",
    x"61E5",
    x"679E",
    x"6CCB",
    x"7165",
    x"7567",
    x"78CA",
    x"7B8A",
    x"7DA5",
    x"7F15",
    x"7FDB",
    x"7FF4",
    x"7F61",
    x"7E22",
    x"7C3A",
    x"79AA",
    x"7675",
    x"72A2",
    x"6E34",
    x"6931",
    x"63A1",
    x"5D8A",
    x"56F6",
    x"4FEC",
    x"4876",
    x"409F",
    x"3871",
    x"2FF7",
    x"273C",
    x"1E4C",
    x"1533",
    x"0BFE",
    x"02B9",
    x"F970",
    x"F030",
    x"E705",
    x"DDFC",
    x"D521",
    x"CC7F",
    x"C423",
    x"BC17",
    x"B467",
    x"AD1D",
    x"A643",
    x"9FE1",
    x"9A01",
    x"94AB",
    x"8FE5",
    x"8BB6",
    x"8824",
    x"8533",
    x"82E8",
    x"8145",
    x"804D",
    x"8001",
    x"8062",
    x"816F",
    x"8326",
    x"8585",
    x"8889",
    x"8C2F",
    x"9070",
    x"9548",
    x"9AAF",
    x"A09F",
    x"A710",
    x"ADF8",
    x"B54F",
    x"BD0B",
    x"C521",
    x"CD86",
    x"D62F",
    x"DF11",
    x"E81E",
    x"F14C",
    x"FA8E",
    x"03D7",
    x"0D1B",
    x"164E",
    x"1F62",
    x"284C",
    x"3100",
    x"3972",
    x"4196",
    x"4962",
    x"50CB",
    x"57C7",
    x"5E4D",
    x"6454",
    x"69D3",
    x"6EC4",
    x"7320",
    x"76E1",
    x"7A01",
    x"7C7D",
    x"7E52",
    x"7F7C",
    x"7FFA",
    x"7FCC",
    x"7EF2",
    x"7D6D",
    x"7B3E",
    x"786A",
    x"74F3",
    x"70DF",
    x"6C33",
    x"66F5",
    x"612C",
    x"5AE0",
    x"541A",
    x"4CE2",
    x"4543",
    x"3D47",
    x"34F8",
    x"2C61",
    x"238F",
    x"1A8D",
    x"1167",
    x"082A",
    x"FEE1",
    x"F59B",
    x"EC62",
    x"E343",
    x"DA4C",
    x"D187",
    x"C901",
    x"C0C5",
    x"B8DE",
    x"B157",
    x"AA39",
    x"A390",
    x"9D63",
    x"97BB",
    x"929F",
    x"8E17",
    x"8A28",
    x"86D8",
    x"842C",
    x"8226",
    x"80CA",
    x"8019",
    x"8014",
    x"80BC",
    x"8210",
    x"840D",
    x"86B1",
    x"89F8",
    x"8DDF",
    x"925F",
    x"9773",
    x"9D14",
    x"A33A",
    x"A9DE",
    x"B0F5",
    x"B877",
    x"C059",
    x"C891",
    x"D113",
    x"D9D5",
    x"E2CB",
    x"EBE7",
    x"F51F",
    x"FE65",
    x"07AE",
    x"10EC",
    x"1A14",
    x"2318",
    x"2BED",
    x"3487",
    x"3CDA",
    x"44DB",
    x"4C7F",
    x"53BC",
    x"5A89",
    x"60DB",
    x"66AB",
    x"6BF0",
    x"70A4",
    x"74C1",
    x"7840",
    x"7B1D",
    x"7D54",
    x"7EE2",
    x"7FC5",
    x"7FFC",
    x"7F87",
    x"7E66",
    x"7C9A",
    x"7A27",
    x"770F",
    x"7356",
    x"6F02",
    x"6A19",
    x"64A0",
    x"5EA1",
    x"5821",
    x"512B",
    x"49C7",
    x"4200",
    x"39E0",
    x"3172",
    x"28C2",
    x"1FDA",
    x"16C8",
    x"0D97",
    x"0453",
    x"FB0A",
    x"F1C8",
    x"E898",
    x"DF88",
    x"D6A4",
    x"CDF8",
    x"C58F",
    x"BD75",
    x"B5B4",
    x"AE58",
    x"A769",
    x"A0F2",
    x"9AFB",
    x"958D",
    x"90AD",
    x"8C64",
    x"88B6",
    x"85A9",
    x"8341",
    x"8181",
    x"806C",
    x"8002",
    x"8045",
    x"8134",
    x"82CE",
    x"8510",
    x"87F8",
    x"8B82",
    x"8FA9",
    x"9467",
    x"99B7",
    x"9F90",
    x"A5EB",
    x"ACBF",
    x"B403",
    x"BBAE",
    x"C3B5",
    x"CC0E",
    x"D4AC",
    x"DD84",
    x"E68C",
    x"EFB5",
    x"F8F4",
    x"023D",
    x"0B83",
    x"14B9",
    x"1DD3",
    x"26C6",
    x"2F84",
    x"3801",
    x"4034",
    x"4810",
    x"4F8B",
    x"569A",
    x"5D35",
    x"6353",
    x"68EA",
    x"6DF4",
    x"726A",
    x"7646",
    x"7983",
    x"7C1C",
    x"7E0D",
    x"7F55",
    x"7FF1",
    x"7FE1",
    x"7F24",
    x"7DBC",
    x"7BAB",
    x"78F3",
    x"7598",
    x"719E",
    x"6D0C",
    x"67E7",
    x"6235",
    x"5BFF",
    x"554E",
    x"4E29",
    x"469B",
    x"3EAE",
    x"366C",
    x"2DE2",
    x"2519",
    x"1C1E",
    x"12FE",
    x"09C3",
    x"007C",
    x"F734",
    x"EDF8",
    x"E4D4",
    x"DBD5",
    x"D306",
    x"CA75",
    x"C22B",
    x"BA34",
    x"B29C",
    x"AB6C",
    x"A4AE",
    x"9E6B",
    x"98AB",
    x"9377",
    x"8ED5",
    x"8ACB",
    x"875F",
    x"8496",
    x"8273",
    x"80FA",
    x"802B",
    x"8009",
    x"8093",
    x"81C9",
    x"83A9",
    x"8630",
    x"895C",
    x"8D27",
    x"918D",
    x"9688",
    x"9C12",
    x"A221",
    x"A8B0",
    x"AFB4",
    x"B724",
    x"BEF6",
    x"C720",
    x"CF96",
    x"D84E",
    x"E13C",
    x"EA52",
    x"F386",
    x"FCCB",
    x"0614",
    x"0F55",
    x"1881",
    x"218C",
    x"2A6A",
    x"330F",
    x"3B6F",
    x"437F",
    x"4B34",
    x"5284",
    x"5965",
    x"5FCD",
    x"65B4",
    x"6B11",
    x"6FDF",
    x"7416",
    x"77B1",
    x"7AAA",
    x"7CFE",
    x"7EA9",
    x"7FAA",
    x"7FFF",
    x"7FA7",
    x"7EA4",
    x"7CF5",
    x"7A9F",
    x"77A3",
    x"7406",
    x"6FCC",
    x"6AFC",
    x"659C",
    x"5FB3",
    x"5949",
    x"5267",
    x"4B15",
    x"435F",
    x"3B4D",
    x"32EC",
    x"2A46",
    x"2167",
    x"185B",
    x"0F2F",
    x"05EE",
    x"FCA5",
    x"F360",
    x"EA2C",
    x"E116",
    x"D82A",
    x"CF73",
    x"C6FD",
    x"BED5",
    x"B704",
    x"AF96",
    x"A894",
    x"A207",
    x"9BFA",
    x"9673",
    x"917A",
    x"8D16",
    x"894D",
    x"8624",
    x"83A0",
    x"81C2",
    x"808F",
    x"8008",
    x"802D",
    x"80FE",
    x"827B",
    x"84A0",
    x"876C",
    x"8ADA",
    x"8EE7",
    x"938B",
    x"98C2",
    x"9E84",
    x"A4C9",
    x"AB89",
    x"B2BB",
    x"BA55",
    x"C24C",
    x"CA97",
    x"D32A",
    x"DBFA",
    x"E4FA",
    x"EE1E",
    x"F75A",
    x"00A2",
    x"09EA",
    x"1324",
    x"1C44",
    x"253E",
    x"2E05",
    x"368F",
    x"3ECF",
    x"46BB",
    x"4E47",
    x"556A",
    x"5C1A",
    x"624E",
    x"67FD",
    x"6D20",
    x"71B0",
    x"75A7",
    x"78FF",
    x"7BB5",
    x"7DC3",
    x"7F28",
    x"7FE2",
    x"7FF0",
    x"7F51",
    x"7E06",
    x"7C12",
    x"7977",
    x"7638",
    x"7259",
    x"6DE1",
    x"68D4",
    x"633A",
    x"5D1B",
    x"567E",
    x"4F6D",
    x"47F0",
    x"4013",
    x"37DF",
    x"2F60",
    x"26A1",
    x"1DAE",
    x"1493",
    x"0B5D",
    x"0217",
    x"F8CE",
    x"EF8F",
    x"E666",
    x"DD5F",
    x"D488",
    x"CBEB",
    x"C394",
    x"BB8E",
    x"B3E5",
    x"ACA2",
    x"A5CF",
    x"9F76",
    x"999F",
    x"9453",
    x"8F97",
    x"8B72",
    x"87EB",
    x"8506",
    x"82C6",
    x"812F",
    x"8042",
    x"8002",
    x"806F",
    x"8187",
    x"834A",
    x"85B5",
    x"88C4",
    x"8C74",
    x"90C0",
    x"95A2",
    x"9B13",
    x"A10C",
    x"A785",
    x"AE75",
    x"B5D4",
    x"BD96",
    x"C5B1",
    x"CE1B",
    x"D6C9",
    x"DFAE",
    x"E8BE",
    x"F1EE",
    x"FB31",
    x"047A",
    x"0DBD",
    x"16EE",
    x"2000",
    x"28E6",
    x"3196",
    x"3A03",
    x"4221",
    x"49E7",
    x"5149",
    x"583D",
    x"5EBA",
    x"64B8",
    x"6A2E",
    x"6F15",
    x"7367",
    x"771D",
    x"7A32",
    x"7CA3",
    x"7E6C",
    x"7F8A",
    x"7FFD",
    x"7FC3",
    x"7EDD",
    x"7D4C",
    x"7B12",
    x"7832",
    x"74B1",
    x"7092",
    x"6BDC",
    x"6694",
    x"60C2",
    x"5A6D",
    x"539F",
    x"4C60",
    x"44BA",
    x"3CB8",
    x"3464",
    x"2BC9",
    x"22F3",
    x"19EE",
    x"10C6",
    x"0788",
    x"FE3F",
    x"F4F9",
    x"EBC1",
    x"E2A5",
    x"D9B1",
    x"D0F0",
    x"C86E",
    x"C038",
    x"B857",
    x"B0D7",
    x"A9C1",
    x"A320",
    x"9CFC",
    x"975D",
    x"924B",
    x"8DCD",
    x"89E9",
    x"86A4",
    x"8403",
    x"8209",
    x"80B8",
    x"8013",
    x"801A",
    x"80CE",
    x"822D",
    x"8436",
    x"86E5",
    x"8A37",
    x"8E29",
    x"92B3",
    x"97D1",
    x"9D7C",
    x"A3AB",
    x"AA56",
    x"B175",
    x"B8FE",
    x"C0E6",
    x"C923",
    x"D1AB",
    x"DA71",
    x"E369",
    x"EC88",
    x"F5C1",
    x"FF08",
    x"0850",
    x"118D",
    x"1AB3",
    x"23B4",
    x"2C85",
    x"351B",
    x"3D68",
    x"4564",
    x"4D01",
    x"5437",
    x"5AFB",
    x"6145",
    x"670B",
    x"6C47",
    x"70F1",
    x"7503",
    x"7877",
    x"7B49",
    x"7D74",
    x"7EF7",
    x"7FCE",
    x"7FFA",
    x"7F78",
    x"7E4C",
    x"7C74",
    x"79F6",
    x"76D3",
    x"730F",
    x"6EB1",
    x"69BE",
    x"643C",
    x"5E33",
    x"57AB",
    x"50AD",
    x"4942",
    x"4175",
    x"394F",
    x"30DC",
    x"2828",
    x"1F3D",
    x"1628",
    x"0CF5",
    x"03B1",
    x"FA68",
    x"F126",
    x"E7F9",
    x"DEEB",
    x"D60B",
    x"CD63",
    x"C4FF",
    x"BCEA",
    x"B530",
    x"ADDB",
    x"A6F4",
    x"A086",
    x"9A98",
    x"9533",
    x"905D",
    x"8C1E",
    x"887C",
    x"857A",
    x"831D",
    x"8169",
    x"805F",
    x"8001",
    x"8050",
    x"814A",
    x"82F0",
    x"853E",
    x"8831",
    x"8BC6",
    x"8FF7",
    x"94C0",
    x"9A19",
    x"9FFB",
    x"A65E",
    x"AD3B",
    x"B486",
    x"BC38",
    x"C445",
    x"CCA2",
    x"D545",
    x"DE21",
    x"E72B",
    x"F056",
    x"F996",
    x"02DF",
    x"0C25",
    x"1559",
    x"1E71",
    x"2760",
    x"301A",
    x"3893",
    x"40C0",
    x"4896",
    x"500A",
    x"5712",
    x"5DA4",
    x"63B9",
    x"6947",
    x"6E47",
    x"72B3",
    x"7684",
    x"79B5",
    x"7C43",
    x"7E29",
    x"7F65",
    x"7FF5",
    x"7FD9",
    x"7F11",
    x"7D9D",
    x"7B80",
    x"78BD",
    x"7557",
    x"7153",
    x"6CB7",
    x"6787",
    x"61CD",
    x"5B8E",
    x"54D4",
    x"4DA8",
    x"4613",
    x"3E20",
    x"35D9",
    x"2D4A",
    x"247D",
    x"1B80",
    x"125D",
    x"0921",
    x"FFDA",
    x"F692",
    x"ED57",
    x"E435",
    x"DB39",
    x"D26E",
    x"C9E1",
    x"C19D",
    x"B9AC",
    x"B21B",
    x"AAF2",
    x"A43C",
    x"9E02",
    x"984C",
    x"9321",
    x"8E89",
    x"8A8A",
    x"8729",
    x"846B",
    x"8254",
    x"80E6",
    x"8023",
    x"800D",
    x"80A3",
    x"81E4",
    x"83D0",
    x"8662",
    x"8999",
    x"8D6F",
    x"91E0",
    x"96E5",
    x"9C77",
    x"A290",
    x"A927",
    x"B032",
    x"B7A9",
    x"BF82",
    x"C7B2",
    x"D02D",
    x"D8E9",
    x"E1D9",
    x"EAF2",
    x"F428",
    x"FD6D",
    x"06B6",
    x"0FF6",
    x"1921",
    x"2229",
    x"2B04",
    x"33A4",
    x"3BFF",
    x"4409",
    x"4BB8",
    x"5300",
    x"59D9",
    x"6038",
    x"6616",
    x"6B6A",
    x"702E",
    x"745A",
    x"77EA",
    x"7AD8",
    x"7D20",
    x"7EC0",
    x"7FB5",
    x"7FFE",
    x"7F9B",
    x"7E8C",
    x"7CD2",
    x"7A70",
    x"7769",
    x"73C1",
    x"6F7D",
    x"6AA3",
    x"6539",
    x"5F47",
    x"58D4",
    x"51EA",
    x"4A91",
    x"42D4",
    x"3ABD",
    x"3257",
    x"29AD",
    x"20CA",
    x"17BC",
    x"0E8D",
    x"054B",
    x"FC02",
    x"F2BE",
    x"E98C",
    x"E079",
    x"D78F",
    x"CEDD",
    x"C66C",
    x"BE49",
    x"B67F",
    x"AF17",
    x"A81D",
    x"A199",
    x"9B95",
    x"9617",
    x"9128",
    x"8CCF",
    x"8911",
    x"85F3",
    x"837A",
    x"81A8",
    x"8081",
    x"8005",
    x"8036",
    x"8113",
    x"829B",
    x"84CC",
    x"87A3",
    x"8B1C",
    x"8F33",
    x"93E2",
    x"9922",
    x"9EED",
    x"A53B",
    x"AC03",
    x"B33C",
    x"BADD",
    x"C2DB",
    x"CB2B",
    x"D3C3",
    x"DC96",
    x"E599",
    x"EEBF",
    x"F7FD",
    x"0145",
    x"0A8C",
    x"13C4",
    x"1CE2",
    x"25D9",
    x"2E9D",
    x"3722",
    x"3F5D",
    x"4742",
    x"4EC8",
    x"55E3",
    x"5C8B",
    x"62B5",
    x"685B",
    x"6D75",
    x"71FA",
    x"75E7",
    x"7934",
    x"7BDE",
    x"7DE1",
    x"7F3B",
    x"7FE9",
    x"7FEA",
    x"7F40",
    x"7DEA",
    x"7BEA",
    x"7943",
    x"75F9",
    x"7210",
    x"6D8D",
    x"6877",
    x"62D3",
    x"5CAB",
    x"5606",
    x"4EED",
    x"4769",
    x"3F86",
    x"374D",
    x"2EC9",
    x"2606",
    x"1D10",
    x"13F3",
    x"0ABB",
    x"0174",
    x"F82C",
    x"EEEE",
    x"E5C7",
    x"DCC3",
    x"D3EF",
    x"CB56",
    x"C304",
    x"BB05",
    x"B362",
    x"AC27",
    x"A55C",
    x"9F0C",
    x"993E",
    x"93FB",
    x"8F49",
    x"8B30",
    x"87B3",
    x"84D9",
    x"82A5",
    x"8119",
    x"8039",
    x"8004",
    x"807D",
    x"81A1",
    x"836F",
    x"85E5",
    x"8900",
    x"8CBB",
    x"9111",
    x"95FD",
    x"9B77",
    x"A179",
    x"A7FB",
    x"AEF3",
    x"B658",
    x"BE21",
    x"C642",
    x"CEB1",
    x"D763",
    x"E04B",
    x"E95E",
    x"F28F",
    x"FBD3",
    x"051C",
    x"0E5F",
    x"178E",
    x"209D",
    x"2980",
    x"322B",
    x"3A93",
    x"42AC",
    x"4A6B",
    x"51C6",
    x"58B2",
    x"5F27",
    x"651C",
    x"6A89",
    x"6F66",
    x"73AD",
    x"7758",
    x"7A62",
    x"7CC7",
    x"7E85",
    x"7F97",
    x"7FFE",
    x"7FB9",
    x"7EC7",
    x"7D2A",
    x"7AE5",
    x"77FA",
    x"746E",
    x"7044",
    x"6B84",
    x"6632",
    x"6057",
    x"59FA",
    x"5324",
    x"4BDE",
    x"4431",
    x"3C29",
    x"33CF",
    x"2B30",
    x"2257",
    x"194F",
    x"1025",
    x"06E5",
    x"FD9D",
    x"F457",
    x"EB21",
    x"E207",
    x"D916",
    x"D059",
    x"C7DC",
    x"BFAB",
    x"B7D0",
    x"B057",
    x"A949",
    x"A2B0",
    x"9C95",
    x"9700",
    x"91F8",
    x"8D84",
    x"89AB",
    x"8671",
    x"83DB",
    x"81EC",
    x"80A7",
    x"800E",
    x"8021",
    x"80E1",
    x"824B",
    x"845F",
    x"871A",
    x"8A77",
    -- nota 02
    x"0000",
    x"09D5",
    x"139A",
    x"1D43",
    x"26BE",
    x"3000",
    x"38F8",
    x"419B",
    x"49DA",
    x"51AA",
    x"58FE",
    x"5FCC",
    x"6608",
    x"6BAB",
    x"70AA",
    x"74FF",
    x"78A3",
    x"7B91",
    x"7DC4",
    x"7F39",
    x"7FED",
    x"7FE0",
    x"7F11",
    x"7D82",
    x"7B36",
    x"782F",
    x"7472",
    x"7005",
    x"6AEF",
    x"6537",
    x"5EE6",
    x"5806",
    x"50A0",
    x"48C1",
    x"4073",
    x"37C4",
    x"2EC0",
    x"2576",
    x"1BF4",
    x"1247",
    x"087E",
    x"FEA8",
    x"F4D5",
    x"EB12",
    x"E16F",
    x"D7FB",
    x"CEC2",
    x"C5D5",
    x"BD3F",
    x"B50E",
    x"AD4F",
    x"A60C",
    x"9F52",
    x"992A",
    x"939D",
    x"8EB4",
    x"8A77",
    x"86EB",
    x"8417",
    x"81FE",
    x"80A3",
    x"8009",
    x"8031",
    x"811A",
    x"82C3",
    x"8529",
    x"8849",
    x"8C1E",
    x"90A2",
    x"95CF",
    x"9B9C",
    x"A202",
    x"A8F5",
    x"B06C",
    x"B85B",
    x"C0B7",
    x"C972",
    x"D280",
    x"DBD3",
    x"E55C",
    x"EF0E",
    x"F8D9",
    x"02AF",
    x"0C81",
    x"1640",
    x"1FDE",
    x"294B",
    x"327A",
    x"3B5D",
    x"43E5",
    x"4C07",
    x"53B6",
    x"5AE7",
    x"618E",
    x"67A1",
    x"6D18",
    x"71EA",
    x"760F",
    x"7982",
    x"7C3D",
    x"7E3D",
    x"7F7D",
    x"7FFD",
    x"7FBB",
    x"7EB7",
    x"7CF4",
    x"7A75",
    x"773C",
    x"734E",
    x"6EB3",
    x"6970",
    x"638D",
    x"5D14",
    x"560E",
    x"4E86",
    x"4687",
    x"3E1E",
    x"3556",
    x"2C3E",
    x"22E3",
    x"1953",
    x"0F9D",
    x"05D0",
    x"FBF9",
    x"F229",
    x"E86D",
    x"DED6",
    x"D570",
    x"CC4B",
    x"C374",
    x"BAF8",
    x"B2E5",
    x"AB47",
    x"A428",
    x"9D95",
    x"9796",
    x"9236",
    x"8D7B",
    x"896E",
    x"8613",
    x"8372",
    x"818C",
    x"8066",
    x"8001",
    x"805D",
    x"817B",
    x"8358",
    x"85F1",
    x"8943",
    x"8D48",
    x"91FB",
    x"9755",
    x"9D4C",
    x"A3D9",
    x"AAF2",
    x"B28B",
    x"BA99",
    x"C310",
    x"CBE3",
    x"D505",
    x"DE68",
    x"E7FE",
    x"F1B8",
    x"FB88",
    x"055E",
    x"0F2D",
    x"18E4",
    x"2276",
    x"2BD3",
    x"34EF",
    x"3DBA",
    x"4628",
    x"4E2C",
    x"55BA",
    x"5CC6",
    x"6345",
    x"692F",
    x"6E79",
    x"731D",
    x"7712",
    x"7A53",
    x"7CDC",
    x"7EA7",
    x"7FB3",
    x"7FFE",
    x"7F87",
    x"7E4F",
    x"7C59",
    x"79A6",
    x"763B",
    x"721E",
    x"6D53",
    x"67E4",
    x"61D7",
    x"5B37",
    x"540C",
    x"4C63",
    x"4446",
    x"3BC1",
    x"32E2",
    x"29B7",
    x"204C",
    x"16B0",
    x"0CF2",
    x"0321",
    x"F94B",
    x"EF7E",
    x"E5CB",
    x"DC40",
    x"D2EA",
    x"C9D9",
    x"C11A",
    x"B8B9",
    x"B0C5",
    x"A948",
    x"A24F",
    x"9BE3",
    x"960F",
    x"90DB",
    x"8C4F",
    x"8871",
    x"8549",
    x"82DA",
    x"8129",
    x"8037",
    x"8007",
    x"8098",
    x"81EA",
    x"83FB",
    x"86C7",
    x"8A4A",
    x"8E80",
    x"9361",
    x"98E6",
    x"9F08",
    x"A5BC",
    x"ACF8",
    x"B4B2",
    x"BCDE",
    x"C570",
    x"CE5A",
    x"D78F",
    x"E101",
    x"EAA2",
    x"F464",
    x"FE37",
    x"080D",
    x"11D6",
    x"1B85",
    x"250A",
    x"2E57",
    x"375E",
    x"4011",
    x"4863",
    x"5048",
    x"57B3",
    x"5E9A",
    x"64F2",
    x"6AB1",
    x"6FCE",
    x"7443",
    x"7808",
    x"7B17",
    x"7D6C",
    x"7F03",
    x"7FDB",
    x"7FF1",
    x"7F45",
    x"7DD9",
    x"7BAF",
    x"78C9",
    x"752D",
    x"70E0",
    x"6BE8",
    x"664D",
    x"6017",
    x"5950",
    x"5201",
    x"4A37",
    x"41FC",
    x"395E",
    x"3069",
    x"272B",
    x"1DB1",
    x"140B",
    x"0A46",
    x"0072",
    x"F69D",
    x"ECD6",
    x"E32C",
    x"D9AE",
    x"D06A",
    x"C76D",
    x"BEC7",
    x"B683",
    x"AEAE",
    x"A754",
    x"A080",
    x"9A3D",
    x"9493",
    x"8F8C",
    x"8B2F",
    x"8783",
    x"848D",
    x"8251",
    x"80D4",
    x"8017",
    x"801B",
    x"80E1",
    x"8268",
    x"84AC",
    x"87AA",
    x"8B5F",
    x"8FC4",
    x"94D3",
    x"9A83",
    x"A0CE",
    x"A7A8",
    x"AF08",
    x"B6E2",
    x"BF2B",
    x"C7D6",
    x"D0D6",
    x"DA1D",
    x"E39E",
    x"ED49",
    x"F711",
    x"00E6",
    x"0ABA",
    x"147E",
    x"1E22",
    x"2799",
    x"30D5",
    x"39C6",
    x"4260",
    x"4A96",
    x"525B",
    x"59A3",
    x"6064",
    x"6692",
    x"6C26",
    x"7117",
    x"755C",
    x"78F0",
    x"7BCC",
    x"7DEE",
    x"7F51",
    x"7FF4",
    x"7FD5",
    x"7EF5",
    x"7D54",
    x"7AF7",
    x"77DF",
    x"7412",
    x"6F95",
    x"6A70",
    x"64AA",
    x"5E4B",
    x"575E",
    x"4FED",
    x"4803",
    x"3FAC",
    x"36F4",
    x"2DEA",
    x"249A",
    x"1B13",
    x"1163",
    x"0798",
    x"FDC2",
    x"F3F0",
    x"EA2F",
    x"E090",
    x"D720",
    x"CDEE",
    x"C508",
    x"BC7B",
    x"B454",
    x"ACA0",
    x"A569",
    x"9EBC",
    x"98A1",
    x"9323",
    x"8E4A",
    x"8A1D",
    x"86A2",
    x"83DE",
    x"81D6",
    x"808D",
    x"8005",
    x"803E",
    x"8139",
    x"82F3",
    x"856A",
    x"889B",
    x"8C81",
    x"9115",
    x"9650",
    x"9C2C",
    x"A29E",
    x"A99E",
    x"B121",
    x"B91A",
    x"C17F",
    x"CA43",
    x"D357",
    x"DCB0",
    x"E63D",
    x"EFF2",
    x"F9BF",
    x"0395",
    x"0D66",
    x"1723",
    x"20BD",
    x"2A25",
    x"334D",
    x"3C28",
    x"44A8",
    x"4CC0",
    x"5464",
    x"5B88",
    x"6222",
    x"6828",
    x"6D90",
    x"7252",
    x"7667",
    x"79CA",
    x"7C74",
    x"7E62",
    x"7F91",
    x"7FFF",
    x"7FAB",
    x"7E96",
    x"7CC2",
    x"7A31",
    x"76E7",
    x"72EA",
    x"6E3E",
    x"68EC",
    x"62FC",
    x"5C75",
    x"5563",
    x"4DD0",
    x"45C7",
    x"3D54",
    x"3485",
    x"2B66",
    x"2206",
    x"1872",
    x"0EB9",
    x"04EA",
    x"FB13",
    x"F144",
    x"E78B",
    x"DDF8",
    x"D497",
    x"CB79",
    x"C2A9",
    x"BA37",
    x"B22E",
    x"AA9B",
    x"A389",
    x"9D02",
    x"9712",
    x"91C0",
    x"8D15",
    x"8918",
    x"85CE",
    x"833D",
    x"8169",
    x"8055",
    x"8001",
    x"8070",
    x"819F",
    x"838D",
    x"8637",
    x"899A",
    x"8DAF",
    x"9272",
    x"97DA",
    x"9DE0",
    x"A47A",
    x"AB9E",
    x"B342",
    x"BB5A",
    x"C3DA",
    x"CCB5",
    x"D5DE",
    x"DF46",
    x"E8E0",
    x"F29D",
    x"FC6E",
    x"0644",
    x"1011",
    x"19C6",
    x"2353",
    x"2CAB",
    x"35C0",
    x"3E83",
    x"46E8",
    x"4EE2",
    x"5664",
    x"5D64",
    x"63D6",
    x"69B1",
    x"6EED",
    x"7381",
    x"7766",
    x"7A96",
    x"7D0E",
    x"7EC8",
    x"7FC2",
    x"7FFB",
    x"7F72",
    x"7E29",
    x"7C21",
    x"795D",
    x"75E2",
    x"71B5",
    x"6CDB",
    x"675D",
    x"6142",
    x"5A95",
    x"535E",
    x"4BAA",
    x"4383",
    x"3AF5",
    x"320F",
    x"28DD",
    x"1F6D",
    x"15CE",
    x"0C0D",
    x"023B",
    x"F865",
    x"EE9A",
    x"E4EA",
    x"DB63",
    x"D213",
    x"C909",
    x"C052",
    x"B7FB",
    x"B011",
    x"A8A0",
    x"A1B3",
    x"9B54",
    x"958E",
    x"9069",
    x"8BED",
    x"8820",
    x"8508",
    x"82AB",
    x"810B",
    x"802B",
    x"800C",
    x"80AF",
    x"8213",
    x"8434",
    x"8711",
    x"8AA5",
    x"8EEB",
    x"93DB",
    x"996F",
    x"9F9E",
    x"A65F",
    x"ADA8",
    x"B56D",
    x"BDA2",
    x"C63D",
    x"CF2E",
    x"D869",
    x"E1E0",
    x"EB85",
    x"F549",
    x"FF1D",
    x"08F2",
    x"12BA",
    x"1C65",
    x"25E6",
    x"2F2D",
    x"382D",
    x"40D8",
    x"4920",
    x"50FA",
    x"585A",
    x"5F34",
    x"657E",
    x"6B2F",
    x"703E",
    x"74A2",
    x"7857",
    x"7B55",
    x"7D99",
    x"7F1F",
    x"7FE5",
    x"7FE9",
    x"7F2C",
    x"7DAE",
    x"7B73",
    x"787C",
    x"74D0",
    x"7073",
    x"6B6B",
    x"65C2",
    x"5F7E",
    x"58AA",
    x"5150",
    x"497B",
    x"4137",
    x"3890",
    x"2F94",
    x"264F",
    x"1CD1",
    x"1327",
    x"0960",
    x"FF8C",
    x"F5B7",
    x"EBF2",
    x"E24C",
    x"D8D3",
    x"CF94",
    x"C69F",
    x"BE01",
    x"B5C7",
    x"ADFD",
    x"A6AE",
    x"9FE7",
    x"99B2",
    x"9417",
    x"8F1F",
    x"8AD2",
    x"8736",
    x"8451",
    x"8227",
    x"80BB",
    x"800F",
    x"8026",
    x"80FD",
    x"8295",
    x"84EA",
    x"87F9",
    x"8BBE",
    x"9033",
    x"9551",
    x"9B10",
    x"A168",
    x"A84F",
    x"AFBA",
    x"B79F",
    x"BFF2",
    x"C8A5",
    x"D1AC",
    x"DAF9",
    x"E47E",
    x"EE2D",
    x"F7F6",
    x"01CC",
    x"0B9F",
    x"1561",
    x"1F02",
    x"2874",
    x"31A9",
    x"3A93",
    x"4324",
    x"4B50",
    x"530A",
    x"5A46",
    x"60FA",
    x"671B",
    x"6CA1",
    x"7182",
    x"75B7",
    x"793A",
    x"7C06",
    x"7E16",
    x"7F68",
    x"7FF9",
    x"7FC8",
    x"7ED7",
    x"7D25",
    x"7AB6",
    x"778E",
    x"73B0",
    x"6F24",
    x"69F0",
    x"641B",
    x"5DAF",
    x"56B6",
    x"4F39",
    x"4744",
    x"3EE4",
    x"3624",
    x"2D13",
    x"23BD",
    x"1A32",
    x"107F",
    x"06B3",
    x"FCDC",
    x"F30B",
    x"E94D",
    x"DFB1",
    x"D647",
    x"CD1B",
    x"C43C",
    x"BBB8",
    x"B39B",
    x"ABF2",
    x"A4C7",
    x"9E27",
    x"981A",
    x"92AB",
    x"8DE1",
    x"89C4",
    x"8659",
    x"83A7",
    x"81B0",
    x"8079",
    x"8002",
    x"804D",
    x"8159",
    x"8325",
    x"85AD",
    x"88EF",
    x"8CE4",
    x"9188",
    x"96D3",
    x"9CBC",
    x"A33C",
    x"AA48",
    x"B1D6",
    x"B9DA",
    x"C248",
    x"CB14",
    x"D42F",
    x"DD8D",
    x"E71F",
    x"F0D6",
    x"FAA5",
    x"047B",
    x"0E4B",
    x"1805",
    x"219B",
    x"2AFE",
    x"3420",
    x"3CF3",
    x"456A",
    x"4D78",
    x"5510",
    x"5C29",
    x"62B5",
    x"68AD",
    x"6E06",
    x"72B9",
    x"76BE",
    x"7A10",
    x"7CA9",
    x"7E86",
    x"7FA3",
    x"7FFF",
    x"7F9A",
    x"7E73",
    x"7C8E",
    x"79EC",
    x"7691",
    x"7284",
    x"6DC9",
    x"6868",
    x"6269",
    x"5BD6",
    x"54B7",
    x"4D18",
    x"4505",
    x"3C8A",
    x"33B3",
    x"2A8D",
    x"2128",
    x"1790",
    x"0DD4",
    x"0404",
    x"FA2D",
    x"F060",
    x"E6AA",
    x"DD1A",
    x"D3BF",
    x"CAA7",
    x"C1E0",
    x"B977",
    x"B178",
    x"A9F0",
    x"A2EA",
    x"9C71",
    x"968F",
    x"914C",
    x"8CB0",
    x"88C3",
    x"858A",
    x"830B",
    x"8148",
    x"8045",
    x"8003",
    x"8083",
    x"81C4",
    x"83C3",
    x"867F",
    x"89F2",
    x"8E17",
    x"92E9",
    x"9860",
    x"9E74",
    x"A51B",
    x"AC4C",
    x"B3FB",
    x"BC1D",
    x"C4A6",
    x"CD89",
    x"D6B7",
    x"E025",
    x"E9C2",
    x"F382",
    x"FD54",
    x"072A",
    x"10F5",
    x"1AA7",
    x"2430",
    x"2D83",
    x"3690",
    x"3F4C",
    x"47A7",
    x"4F96",
    x"570D",
    x"5E00",
    x"6465",
    x"6A32",
    x"6F5F",
    x"73E3",
    x"77B8",
    x"7AD8",
    x"7D3E",
    x"7EE6",
    x"7FCF",
    x"7FF6",
    x"7F5C",
    x"7E02",
    x"7BE8",
    x"7914",
    x"7588",
    x"714A",
    x"6C61",
    x"66D5",
    x"60AC",
    x"59F2",
    x"52AF",
    x"4AF0",
    x"42BF",
    x"3A29",
    x"313B",
    x"2803",
    x"1E8E",
    x"14EB",
    x"0B28",
    x"0155",
    x"F77F",
    x"EDB7",
    x"E40A",
    x"DA87",
    x"D13D",
    x"C839",
    x"BF8B",
    x"B73D",
    x"AF5E",
    x"A7F8",
    x"A118",
    x"9AC7",
    x"950F",
    x"8FF9",
    x"8B8D",
    x"87D0",
    x"84C9",
    x"827D",
    x"80EF",
    x"8020",
    x"8013",
    x"80C8",
    x"823D",
    x"8470",
    x"875E",
    x"8B02",
    x"8F57",
    x"9457",
    x"99FA",
    x"A036",
    x"A704",
    x"AE58",
    x"B628",
    x"BE68",
    x"C70A",
    x"D003",
    x"D944",
    x"E2C0",
    x"EC68",
    x"F62E",
    x"0003",
    x"09D8",
    x"139D",
    x"1D45",
    x"26C1",
    x"3002",
    x"38FB",
    x"419D",
    x"49DD",
    x"51AC",
    x"5900",
    x"5FCD",
    x"660A",
    x"6BAC",
    x"70AB",
    x"7500",
    x"78A4",
    x"7B92",
    x"7DC5",
    x"7F39",
    x"7FED",
    x"7FE0",
    x"7F11",
    x"7D82",
    x"7B35",
    x"782E",
    x"7471",
    x"7004",
    x"6AEE",
    x"6536",
    x"5EE4",
    x"5804",
    x"509E",
    x"48BE",
    x"4070",
    x"37C1",
    x"2EBE",
    x"2574",
    x"1BF1",
    x"1244",
    x"087B",
    x"FEA5",
    x"F4D2",
    x"EB0F",
    x"E16C",
    x"D7F8",
    x"CEC0",
    x"C5D2",
    x"BD3C",
    x"B50C",
    x"AD4C",
    x"A60A",
    x"9F50",
    x"9928",
    x"939C",
    x"8EB3",
    x"8A76",
    x"86EB",
    x"8416",
    x"81FD",
    x"80A3",
    x"8009",
    x"8031",
    x"811A",
    x"82C3",
    x"852A",
    x"884A",
    x"8C1F",
    x"90A4",
    x"95D1",
    x"9B9E",
    x"A204",
    x"A8F7",
    x"B06E",
    x"B85E",
    x"C0B9",
    x"C975",
    x"D283",
    x"DBD6",
    x"E55F",
    x"EF11",
    x"F8DC",
    x"02B2",
    x"0C84",
    x"1643",
    x"1FE1",
    x"294E",
    x"327D",
    x"3B5F",
    x"43E8",
    x"4C0A",
    x"53B9",
    x"5AE9",
    x"6190",
    x"67A3",
    x"6D1A",
    x"71EB",
    x"7610",
    x"7983",
    x"7C3E",
    x"7E3D",
    x"7F7D",
    x"7FFD",
    x"7FBA",
    x"7EB7",
    x"7CF4",
    x"7A74",
    x"773B",
    x"734D",
    x"6EB1",
    x"696E",
    x"638B",
    x"5D12",
    x"560C",
    x"4E84",
    x"4685",
    x"3E1B",
    x"3554",
    x"2C3B",
    x"22E0",
    x"1951",
    x"0F9A",
    x"05CD",
    x"FBF6",
    x"F226",
    -- nota 03
    x"0000",
    x"0A6A",
    x"14C2",
    x"1EF8",
    x"28F8",
    x"32B3",
    x"3C18",
    x"4517",
    x"4DA1",
    x"55A6",
    x"5D1B",
    x"63F1",
    x"6A1E",
    x"6F97",
    x"7452",
    x"7848",
    x"7B71",
    x"7DC9",
    x"7F4C",
    x"7FF6",
    x"7FC7",
    x"7EC0",
    x"7CE1",
    x"7A2E",
    x"76AC",
    x"7260",
    x"6D52",
    x"678A",
    x"6113",
    x"59F7",
    x"5242",
    x"4A02",
    x"4144",
    x"3817",
    x"2E8B",
    x"24B0",
    x"1A97",
    x"1050",
    x"05EE",
    x"FB82",
    x"F11E",
    x"E6D2",
    x"DCB2",
    x"D2CD",
    x"C935",
    x"BFFA",
    x"B72C",
    x"AED9",
    x"A711",
    x"9FDF",
    x"9950",
    x"9370",
    x"8E48",
    x"89E1",
    x"8642",
    x"8372",
    x"8176",
    x"8050",
    x"8003",
    x"8090",
    x"81F4",
    x"842F",
    x"873C",
    x"8B16",
    x"8FB6",
    x"9515",
    x"9B2A",
    x"A1E9",
    x"A949",
    x"B13B",
    x"B9B4",
    x"C2A3",
    x"CBFB",
    x"D5AB",
    x"DFA3",
    x"E9D2",
    x"F427",
    x"FE8F",
    x"08FA",
    x"1356",
    x"1D91",
    x"279A",
    x"3160",
    x"3AD1",
    x"43DF",
    x"4C7A",
    x"5493",
    x"5C1C",
    x"6309",
    x"694E",
    x"6EE0",
    x"73B6",
    x"77C8",
    x"7B0E",
    x"7D83",
    x"7F23",
    x"7FEC",
    x"7FDB",
    x"7EF1",
    x"7D30",
    x"7A9A",
    x"7734",
    x"7304",
    x"6E10",
    x"6862",
    x"6202",
    x"5AFC",
    x"535C",
    x"4B2E",
    x"4280",
    x"3962",
    x"2FE2",
    x"2611",
    x"1BFF",
    x"11BE",
    x"075F",
    x"FCF3",
    x"F28C",
    x"E83C",
    x"DE15",
    x"D427",
    x"CA83",
    x"C13B",
    x"B85C",
    x"AFF8",
    x"A81B",
    x"A0D4",
    x"9A2E",
    x"9435",
    x"8EF3",
    x"8A70",
    x"86B6",
    x"83C9",
    x"81AF",
    x"806C",
    x"8001",
    x"806F",
    x"81B6",
    x"83D4",
    x"86C4",
    x"8A82",
    x"8F07",
    x"944C",
    x"9A48",
    x"A0F1",
    x"A83B",
    x"B01A",
    x"B881",
    x"C161",
    x"CAAB",
    x"D450",
    x"DE3F",
    x"E867",
    x"F2B8",
    x"FD1E",
    x"078A",
    x"11E9",
    x"1C2A",
    x"263B",
    x"300B",
    x"3989",
    x"42A6",
    x"4B51",
    x"537D",
    x"5B1B",
    x"621E",
    x"687B",
    x"6E26",
    x"7317",
    x"7744",
    x"7AA6",
    x"7D39",
    x"7EF7",
    x"7FDD",
    x"7FEA",
    x"7F1E",
    x"7D7A",
    x"7B02",
    x"77B8",
    x"73A3",
    x"6ECA",
    x"6935",
    x"62EE",
    x"5BFE",
    x"5472",
    x"4C57",
    x"43BA",
    x"3AAB",
    x"3137",
    x"2770",
    x"1D67",
    x"132B",
    x"08CF",
    x"FE63",
    x"F3FB",
    x"E9A7",
    x"DF79",
    x"D582",
    x"CBD3",
    x"C27D",
    x"B98F",
    x"B119",
    x"A929",
    x"A1CC",
    x"9B0F",
    x"94FD",
    x"8FA1",
    x"8B04",
    x"872E",
    x"8424",
    x"81ED",
    x"808C",
    x"8003",
    x"8053",
    x"817C",
    x"837C",
    x"8650",
    x"89F1",
    x"8E5C",
    x"9387",
    x"996A",
    x"9FFC",
    x"A730",
    x"AEFB",
    x"B750",
    x"C020",
    x"C95D",
    x"D2F6",
    x"DCDC",
    x"E6FD",
    x"F149",
    x"FBAE",
    x"061A",
    x"107C",
    x"1AC2",
    x"24DA",
    x"2EB4",
    x"383F",
    x"416A",
    x"4A26",
    x"5264",
    x"5A16",
    x"6130",
    x"67A4",
    x"6D69",
    x"7273",
    x"76BC",
    x"7A3B",
    x"7CEA",
    x"7EC6",
    x"7FCA",
    x"7FF5",
    x"7F47",
    x"7DC1",
    x"7B66",
    x"7839",
    x"7440",
    x"6F81",
    x"6A06",
    x"63D6",
    x"5CFD",
    x"5586",
    x"4D7E",
    x"44F2",
    x"3BF1",
    x"328B",
    x"28CF",
    x"1ECD",
    x"1497",
    x"0A3E",
    x"FFD4",
    x"F56A",
    x"EB12",
    x"E0DE",
    x"D6DE",
    x"CD25",
    x"C3C1",
    x"BAC4",
    x"B23D",
    x"AA39",
    x"A2C7",
    x"9BF3",
    x"95C9",
    x"9054",
    x"8B9C",
    x"87A9",
    x"8483",
    x"822F",
    x"80B0",
    x"8009",
    x"803B",
    x"8146",
    x"8329",
    x"85DF",
    x"8965",
    x"8DB4",
    x"92C5",
    x"988F",
    x"9F09",
    x"A628",
    x"ADDF",
    x"B622",
    x"BEE2",
    x"C810",
    x"D19D",
    x"DB7A",
    x"E594",
    x"EFDB",
    x"FA3D",
    x"04AA",
    x"0F0E",
    x"1959",
    x"2378",
    x"2D5C",
    x"36F2",
    x"402C",
    x"48F8",
    x"5148",
    x"590F",
    x"603E",
    x"66CA",
    x"6CA8",
    x"71CC",
    x"7630",
    x"79CB",
    x"7C98",
    x"7E91",
    x"7FB3",
    x"7FFC",
    x"7F6C",
    x"7E04",
    x"7BC6",
    x"78B5",
    x"74D8",
    x"7035",
    x"6AD3",
    x"64BB",
    x"5DF9",
    x"5697",
    x"4EA2",
    x"4628",
    x"3D36",
    x"33DD",
    x"2A2B",
    x"2033",
    x"1603",
    x"0BAE",
    x"0145",
    x"F6DA",
    x"EC7F",
    x"E244",
    x"D83C",
    x"CE78",
    x"C508",
    x"BBFC",
    x"B363",
    x"AB4C",
    x"A3C5",
    x"9CDB",
    x"9699",
    x"910A",
    x"8C37",
    x"8829",
    x"84E6",
    x"8274",
    x"80D8",
    x"8013",
    x"8027",
    x"8115",
    x"82DA",
    x"8573",
    x"88DC",
    x"8D10",
    x"9206",
    x"97B8",
    x"9E1A",
    x"A523",
    x"ACC6",
    x"B4F6",
    x"BDA5",
    x"C6C5",
    x"D047",
    x"DA19",
    x"E42B",
    x"EE6D",
    x"F8CD",
    x"0339",
    x"0D9F",
    x"17EF",
    x"2215",
    x"2C02",
    x"35A4",
    x"3EEC",
    x"47C8",
    x"502A",
    x"5805",
    x"5F4A",
    x"65ED",
    x"6BE3",
    x"7122",
    x"75A1",
    x"7958",
    x"7C41",
    x"7E58",
    x"7F98",
    x"7FFF",
    x"7F8D",
    x"7E42",
    x"7C22",
    x"792E",
    x"756D",
    x"70E4",
    x"6B9C",
    x"659D",
    x"5EF2",
    x"57A5",
    x"4FC4",
    x"475B",
    x"3E79",
    x"352D",
    x"2B87",
    x"2197",
    x"176E",
    x"0D1D",
    x"02B6",
    x"F84A",
    x"EDEB",
    x"E3AB",
    x"D99C",
    x"CFCD",
    x"C650",
    x"BD35",
    x"B48B",
    x"AC62",
    x"A4C6",
    x"9DC6",
    x"976C",
    x"91C3",
    x"8CD6",
    x"88AC",
    x"854D",
    x"82BE",
    x"8104",
    x"8021",
    x"8018",
    x"80E7",
    x"828E",
    x"850A",
    x"8857",
    x"8C6F",
    x"914B",
    x"96E4",
    x"9D2E",
    x"A420",
    x"ABAF",
    x"B3CC",
    x"BC6B",
    x"C57C",
    x"CEF1",
    x"D8B9",
    x"E2C4",
    x"ED00",
    x"F75D",
    x"01C8",
    x"0C31",
    x"1684",
    x"20B1",
    x"2AA7",
    x"3455",
    x"3DA9",
    x"4695",
    x"4F09",
    x"56F7",
    x"5E52",
    x"650C",
    x"6B1B",
    x"7074",
    x"750D",
    x"78E1",
    x"7BE7",
    x"7E1B",
    x"7F78",
    x"7FFE",
    x"7FAA",
    x"7E7D",
    x"7C7A",
    x"79A3",
    x"75FE",
    x"7190",
    x"6C62",
    x"667C",
    x"5FE7",
    x"58B0",
    x"50E3",
    x"488C",
    x"3FBA",
    x"367C",
    x"2CE1",
    x"22FA",
    x"18D8",
    x"0E8C",
    x"0426",
    x"F9BA",
    x"EF59",
    x"E513",
    x"DAFC",
    x"D123",
    x"C79A",
    x"BE71",
    x"B5B7",
    x"AD7B",
    x"A5CB",
    x"9EB4",
    x"9842",
    x"9281",
    x"8D79",
    x"8934",
    x"85B8",
    x"830C",
    x"8134",
    x"8034",
    x"800C",
    x"80BD",
    x"8247",
    x"84A6",
    x"87D6",
    x"8BD3",
    x"9094",
    x"9613",
    x"9C45",
    x"A321",
    x"AA9B",
    x"B2A5",
    x"BB33",
    x"C435",
    x"CD9D",
    x"D75B",
    x"E15D",
    x"EB94",
    x"F5ED",
    x"0057",
    x"0AC1",
    x"1519",
    x"1F4C",
    x"294B",
    x"3303",
    x"3C65",
    x"4561",
    x"4DE6",
    x"55E7",
    x"5D57",
    x"6428",
    x"6A4F",
    x"6FC2",
    x"7476",
    x"7866",
    x"7B88",
    x"7DD9",
    x"7F55",
    x"7FF8",
    x"7FC2",
    x"7EB3",
    x"7CCD",
    x"7A14",
    x"768B",
    x"7238",
    x"6D24",
    x"6757",
    x"60DA",
    x"59B9",
    x"51FF",
    x"49BB",
    x"40F9",
    x"37C9",
    x"2E3A",
    x"245C",
    x"1A41",
    x"0FFA",
    x"0597",
    x"FB2B",
    x"F0C7",
    x"E67C",
    x"DC5E",
    x"D27B",
    x"C8E6",
    x"BFAE",
    x"B6E4",
    x"AE96",
    x"A6D2",
    x"9FA5",
    x"991C",
    x"9341",
    x"8E20",
    x"89BF",
    x"8627",
    x"835E",
    x"8169",
    x"804A",
    x"8004",
    x"8098",
    x"8204",
    x"8446",
    x"8759",
    x"8B3A",
    x"8FE0",
    x"9546",
    x"9B60",
    x"A225",
    x"A989",
    x"B180",
    x"B9FD",
    x"C2F0",
    x"CC4B",
    x"D5FE",
    x"DFF8",
    x"EA28",
    x"F47E",
    x"FEE7",
    x"0952",
    x"13AD",
    x"1DE6",
    x"27ED",
    x"31B0",
    x"3B1F",
    x"442A",
    x"4CC0",
    x"54D5",
    x"5C59",
    x"6341",
    x"6980",
    x"6F0C",
    x"73DC",
    x"77E6",
    x"7B26",
    x"7D94",
    x"7F2D",
    x"7FEE",
    x"7FD7",
    x"7EE6",
    x"7D1D",
    x"7A81",
    x"7714",
    x"72DD",
    x"6DE3",
    x"682F",
    x"61CA",
    x"5ABE",
    x"5319",
    x"4AE7",
    x"4235",
    x"3914",
    x"2F91",
    x"25BD",
    x"1BAA",
    x"1167",
    x"0707",
    x"FC9B",
    x"F235",
    x"E7E6",
    x"DDC0",
    x"D3D5",
    x"CA34",
    x"C0EE",
    x"B814",
    x"AFB4",
    x"A7DC",
    x"A099",
    x"99F9",
    x"9406",
    x"8ECA",
    x"8A4E",
    x"869A",
    x"83B4",
    x"81A1",
    x"8065",
    x"8001",
    x"8077",
    x"81C5",
    x"83E9",
    x"86E0",
    x"8AA5",
    x"8F30",
    x"947C",
    x"9A7E",
    x"A12C",
    x"A87B",
    x"B05E",
    x"B8C9",
    x"C1AD",
    x"CAFB",
    x"D4A2",
    x"DE93",
    x"E8BD",
    x"F30F",
    x"FD76",
    x"07E2",
    x"1240",
    x"1C7F",
    x"268E",
    x"305C",
    x"39D7",
    x"42F0",
    x"4B98",
    x"53BF",
    x"5B58",
    x"6256",
    x"68AD",
    x"6E53",
    x"733D",
    x"7763",
    x"7ABF",
    x"7D4B",
    x"7F02",
    x"7FE1",
    x"7FE7",
    x"7F14",
    x"7D69",
    x"7AE9",
    x"7799",
    x"737E",
    x"6E9F",
    x"6903",
    x"62B6",
    x"5BC1",
    x"5430",
    x"4C11",
    x"4370",
    x"3A5D",
    x"30E6",
    x"271D",
    x"1D11",
    x"12D4",
    x"0877",
    x"FE0C",
    x"F3A4",
    x"E951",
    x"DF24",
    x"D52F",
    x"CB83",
    x"C230",
    x"B946",
    x"B0D4",
    x"A8E8",
    x"A191",
    x"9AD9",
    x"94CD",
    x"8F78",
    x"8AE1",
    x"8711",
    x"840E",
    x"81DE",
    x"8084",
    x"8002",
    x"805A",
    x"818A",
    x"8391",
    x"866B",
    x"8A13",
    x"8E84",
    x"93B5",
    x"999F",
    x"A036",
    x"A76F",
    x"AF3F",
    x"B798",
    x"C06C",
    x"C9AC",
    x"D348",
    x"DD30",
    x"E753",
    x"F1A0",
    x"FC05",
    x"0671",
    x"10D3",
    x"1B17",
    x"252E",
    x"2F05",
    x"388D",
    x"41B5",
    x"4A6D",
    x"52A7",
    x"5A54",
    x"6169",
    x"67D7",
    x"6D96",
    x"729B",
    x"76DD",
    x"7A55",
    x"7CFD",
    x"7ED2",
    x"7FCF",
    x"7FF3",
    x"7F3E",
    x"7DB1",
    x"7B4E",
    x"781B",
    x"741B",
    x"6F56",
    x"69D5",
    x"639F",
    x"5CC1",
    x"5545",
    x"4D38",
    x"44A8",
    x"3BA4",
    x"323A",
    x"287C",
    x"1E78",
    x"1441",
    x"09E7",
    x"FF7D",
    x"F513",
    x"EABC",
    x"E089",
    x"D68C",
    x"CCD5",
    x"C374",
    x"BA7B",
    x"B1F7",
    x"A9F8",
    x"A28B",
    x"9BBD",
    x"9599",
    x"9029",
    x"8B77",
    x"878C",
    x"846C",
    x"821F",
    x"80A7",
    x"8007",
    x"8041",
    x"8153",
    x"833C",
    x"85FA",
    x"8986",
    x"8DDB",
    x"92F3",
    x"98C3",
    x"9F42",
    x"A666",
    x"AE22",
    x"B669",
    x"BF2D",
    x"C85F",
    x"D1EF",
    x"DBCE",
    x"E5EA",
    x"F032",
    x"FA95",
    x"0501",
    x"0F65",
    x"19AE",
    x"23CC",
    x"2DAE",
    x"3741",
    x"4077",
    x"4940",
    x"518C",
    x"594E",
    x"6078",
    x"66FE",
    x"6CD6",
    x"71F4",
    x"7652",
    x"79E6",
    x"7CAC",
    x"7E9E",
    x"7FB9",
    x"7FFB",
    x"7F64",
    x"7DF4",
    x"7BAF",
    x"7898",
    x"74B4",
    x"700A",
    x"6AA2",
    x"6485",
    x"5DBD",
    x"5656",
    x"4E5D",
    x"45DE",
    x"3CE9",
    x"338D",
    x"29D9",
    x"1FDE",
    x"15AD",
    x"0B57",
    x"00EE",
    x"F683",
    x"EC28",
    x"E1EF",
    x"D7E9",
    x"CE27",
    x"C4BA",
    x"BBB1",
    x"B31D",
    x"AB0B",
    x"A389",
    x"9CA4",
    x"9667",
    x"90DE",
    x"8C12",
    x"880A",
    x"84CE",
    x"8263",
    x"80CE",
    x"8010",
    x"802C",
    x"8120",
    x"82EC",
    x"858C",
    x"88FC",
    x"8D36",
    x"9233",
    x"97EB",
    x"9E53",
    x"A560",
    x"AD08",
    x"B53D",
    x"BDF0",
    x"C714",
    x"D098",
    x"DA6C",
    x"E481",
    x"EEC4",
    x"F924",
    x"0390",
    x"0DF6",
    x"1845",
    x"226A",
    x"2C54",
    x"35F4",
    x"3F38",
    x"4810",
    x"506E",
    x"5844",
    x"5F84",
    x"6622",
    x"6C12",
    x"714B",
    x"75C3",
    x"7974",
    x"7C56",
    x"7E66",
    x"7F9E",
    x"7FFF",
    x"7F86",
    x"7E34",
    x"7C0C",
    x"7912",
    x"754A",
    x"70BB",
    x"6B6D",
    x"6568",
    x"5EB7",
    x"5765",
    x"4F7F",
    x"4712",
    x"3E2D",
    x"34DE",
    x"2B35",
    x"2142",
    x"1718",
    x"0CC6",
    x"025E",
    x"F7F3",
    x"ED95",
    x"E356",
    x"D948",
    x"CF7C",
    x"C602",
    x"BCEA",
    x"B445",
    x"AC20",
    x"A489",
    x"9D8E",
    x"9739",
    x"9197",
    x"8CB0",
    x"888D",
    x"8534",
    x"82AC",
    x"80F9",
    x"801D",
    x"801B",
    x"80F1",
    x"82A0",
    x"8523",
    x"8876",
    x"8C95",
    x"9177",
    x"9716",
    x"9D66",
    x"A45D",
    x"ABF1",
    x"B412",
    x"BCB5",
    x"C5CA",
    x"CF42",
    x"D90D",
    x"E319",
    x"ED57",
    x"F7B4",
    x"0220",
    x"0C88",
    x"16DA",
    x"2106",
    x"2AFA",
    x"34A5",
    x"3DF6",
    x"46DE",
    x"4F4E",
    x"5738",
    x"5E8D",
    x"6542",
    x"6B4A",
    x"709D",
    x"7531",
    x"78FD",
    x"7BFD",
    x"7E29",
    x"7F80",
    x"7FFE",
    x"7FA3",
    -- nota 04
    x"0000",
    x"0B08",
    x"15FB",
    x"20C5",
    x"2B4F",
    x"3588",
    x"3F5A",
    x"48B4",
    x"5183",
    x"59B7",
    x"6140",
    x"680F",
    x"6E19",
    x"7350",
    x"77AC",
    x"7B24",
    x"7DB1",
    x"7F4F",
    x"7FFA",
    x"7FB1",
    x"7E75",
    x"7C49",
    x"792F",
    x"752E",
    x"704F",
    x"6A99",
    x"6418",
    x"5CD8",
    x"54E8",
    x"4C56",
    x"4332",
    x"398E",
    x"2F7D",
    x"2511",
    x"1A5E",
    x"0F7A",
    x"0477",
    x"F96D",
    x"EE6F",
    x"E392",
    x"D8EB",
    x"CE8F",
    x"C491",
    x"BB05",
    x"B1FB",
    x"A987",
    x"A1B7",
    x"9A9B",
    x"9440",
    x"8EB2",
    x"89FC",
    x"8627",
    x"833B",
    x"813B",
    x"802E",
    x"8014",
    x"80EE",
    x"82B9",
    x"8574",
    x"8918",
    x"8D9E",
    x"92FF",
    x"992F",
    x"A023",
    x"A7CE",
    x"B021",
    x"B90B",
    x"C27E",
    x"CC65",
    x"D6AE",
    x"E147",
    x"EC1A",
    x"F713",
    x"021C",
    x"0D22",
    x"180F",
    x"22CE",
    x"2D4A",
    x"3771",
    x"412D",
    x"4A6E",
    x"5321",
    x"5B35",
    x"629C",
    x"6946",
    x"6F28",
    x"7437",
    x"7867",
    x"7BB3",
    x"7E13",
    x"7F82",
    x"7FFF",
    x"7F88",
    x"7E1E",
    x"7BC3",
    x"787D",
    x"7451",
    x"6F47",
    x"696A",
    x"62C4",
    x"5B61",
    x"5350",
    x"4AA1",
    x"4164",
    x"37A9",
    x"2D85",
    x"230A",
    x"184D",
    x"0D61",
    x"025B",
    x"F751",
    x"EC58",
    x"E184",
    x"D6EA",
    x"CC9F",
    x"C2B5",
    x"B940",
    x"B052",
    x"A7FB",
    x"A04D",
    x"9955",
    x"9320",
    x"8DBB",
    x"892F",
    x"8586",
    x"82C6",
    x"80F5",
    x"8016",
    x"802B",
    x"8133",
    x"832D",
    x"8614",
    x"89E4",
    x"8E95",
    x"941E",
    x"9A74",
    x"A18C",
    x"A958",
    x"B1CA",
    x"BAD0",
    x"C45A",
    x"CE55",
    x"D8AF",
    x"E354",
    x"EE30",
    x"F92E",
    x"0439",
    x"0F3B",
    x"1A21",
    x"24D5",
    x"2F42",
    x"3956",
    x"42FC",
    x"4C23",
    x"54B9",
    x"5CAD",
    x"63F1",
    x"6A76",
    x"7030",
    x"7515",
    x"791B",
    x"7C39",
    x"7E6C",
    x"7FAD",
    x"7FFB",
    x"7F55",
    x"7DBD",
    x"7B35",
    x"77C2",
    x"736B",
    x"6E39",
    x"6834",
    x"6168",
    x"59E4",
    x"51B3",
    x"48E8",
    x"3F91",
    x"35C1",
    x"2B8B",
    x"2101",
    x"1639",
    x"0B47",
    x"003F",
    x"F537",
    x"EA43",
    x"DF78",
    x"D4EC",
    x"CAB1",
    x"C0DD",
    x"B780",
    x"AEAE",
    x"A676",
    x"9EE9",
    x"9816",
    x"9208",
    x"8CCB",
    x"886A",
    x"84ED",
    x"825B",
    x"80B8",
    x"8007",
    x"804A",
    x"8181",
    x"83A8",
    x"86BD",
    x"8AB8",
    x"8F93",
    x"9544",
    x"9BC1",
    x"A2FC",
    x"AAE9",
    x"B378",
    x"BC99",
    x"C63A",
    x"D049",
    x"DAB3",
    x"E564",
    x"F048",
    x"FB4A",
    x"0654",
    x"1153",
    x"1C31",
    x"26D9",
    x"3137",
    x"3B37",
    x"44C6",
    x"4DD3",
    x"564B",
    x"5E1E",
    x"653F",
    x"6B9E",
    x"7131",
    x"75EB",
    x"79C5",
    x"7CB7",
    x"7EBC",
    x"7FCF",
    x"7FEE",
    x"7F1A",
    x"7D53",
    x"7A9E",
    x"76FF",
    x"727E",
    x"6D22",
    x"66F6",
    x"6007",
    x"5860",
    x"5011",
    x"4729",
    x"3DBA",
    x"33D5",
    x"298D",
    x"1EF6",
    x"1424",
    x"092C",
    x"FE23",
    x"F31D",
    x"E82F",
    x"DD6F",
    x"D2F0",
    x"C8C8",
    x"BF09",
    x"B5C5",
    x"AD0F",
    x"A4F7",
    x"9D8D",
    x"96DE",
    x"90F7",
    x"8BE4",
    x"87AE",
    x"845D",
    x"81F8",
    x"8083",
    x"8001",
    x"8073",
    x"81D8",
    x"842D",
    x"876E",
    x"8B95",
    x"9099",
    x"9672",
    x"9D14",
    x"A473",
    x"AC80",
    x"B52C",
    x"BE66",
    x"C81E",
    x"D240",
    x"DCB9",
    x"E775",
    x"F261",
    x"FD66",
    x"0870",
    x"136A",
    x"1E3F",
    x"28DA",
    x"3328",
    x"3D14",
    x"468C",
    x"4F7D",
    x"57D7",
    x"5F89",
    x"6686",
    x"6CBF",
    x"7229",
    x"76B9",
    x"7A68",
    x"7D2D",
    x"7F03",
    x"7FE8",
    x"7FD8",
    x"7ED6",
    x"7CE1",
    x"79FF",
    x"7634",
    x"7188",
    x"6C04",
    x"65B2",
    x"5E9E",
    x"56D6",
    x"4E68",
    x"4565",
    x"3BDE",
    x"31E5",
    x"278D",
    x"1CE9",
    x"120E",
    x"0711",
    x"FC06",
    x"F103",
    x"E61D",
    x"DB68",
    x"D0F8",
    x"C6E2",
    x"BD39",
    x"B410",
    x"AB77",
    x"A37F",
    x"9C37",
    x"95AD",
    x"8FEE",
    x"8B05",
    x"86FA",
    x"83D6",
    x"819E",
    x"8058",
    x"8004",
    x"80A4",
    x"8237",
    x"84BA",
    x"8828",
    x"8C79",
    x"91A7",
    x"97A8",
    x"9E6F",
    x"A5F0",
    x"AE1C",
    x"B6E5",
    x"C039",
    x"CA06",
    x"D43A",
    x"DEC2",
    x"E989",
    x"F47A",
    x"FF82",
    x"0A8B",
    x"157F",
    x"204B",
    x"2AD9",
    x"3515",
    x"3EED",
    x"484C",
    x"5122",
    x"595D",
    x"60EE",
    x"67C6",
    x"6DD8",
    x"7319",
    x"777F",
    x"7B01",
    x"7D99",
    x"7F42",
    x"7FF8",
    x"7FBA",
    x"7E89",
    x"7C66",
    x"7957",
    x"7561",
    x"708B",
    x"6ADE",
    x"6466",
    x"5D2F",
    x"5546",
    x"4CBA",
    x"439D",
    x"39FE",
    x"2FF2",
    x"2589",
    x"1ADA",
    x"0FF7",
    x"04F5",
    x"F9EA",
    x"EEEB",
    x"E40D",
    x"D963",
    x"CF03",
    x"C501",
    x"BB6F",
    x"B25F",
    x"A9E4",
    x"A20C",
    x"9AE8",
    x"9484",
    x"8EED",
    x"8A2D",
    x"864E",
    x"8357",
    x"814D",
    x"8035",
    x"8010",
    x"80DF",
    x"82A0",
    x"8550",
    x"88EA",
    x"8D66",
    x"92BD",
    x"98E4",
    x"9FD0",
    x"A773",
    x"AFBE",
    x"B8A3",
    x"C20F",
    x"CBF2",
    x"D637",
    x"E0CD",
    x"EB9D",
    x"F695",
    x"019E",
    x"0CA5",
    x"1793",
    x"2255",
    x"2CD5",
    x"36FF",
    x"40C1",
    x"4A07",
    x"52C1",
    x"5ADC",
    x"624B",
    x"68FE",
    x"6EEA",
    x"7402",
    x"783D",
    x"7B92",
    x"7DFD",
    x"7F77",
    x"7FFF",
    x"7F92",
    x"7E33",
    x"7BE3",
    x"78A7",
    x"7485",
    x"6F85",
    x"69B1",
    x"6314",
    x"5BB9",
    x"53B0",
    x"4B07",
    x"41D0",
    x"381B",
    x"2DFB",
    x"2383",
    x"18C8",
    x"0DDE",
    x"02D9",
    x"F7CF",
    x"ECD4",
    x"E1FE",
    x"D761",
    x"CD12",
    x"C323",
    x"B9A9",
    x"B0B4",
    x"A857",
    x"A0A1",
    x"99A0",
    x"9362",
    x"8DF4",
    x"895E",
    x"85AB",
    x"82E1",
    x"8105",
    x"801B",
    x"8025",
    x"8122",
    x"8311",
    x"85EE",
    x"89B4",
    x"8E5B",
    x"93DA",
    x"9A28",
    x"A138",
    x"A8FC",
    x"B166",
    x"BA66",
    x"C3EA",
    x"CDE1",
    x"D838",
    x"E2DA",
    x"EDB3",
    x"F8B0",
    x"03BB",
    x"0EBE",
    x"19A5",
    x"245C",
    x"2ECD",
    x"38E5",
    x"4291",
    x"4BBE",
    x"545A",
    x"5C56",
    x"63A2",
    x"6A30",
    x"6FF3",
    x"74E2",
    x"78F2",
    x"7C1B",
    x"7E58",
    x"7FA4",
    x"7FFD",
    x"7F62",
    x"7DD4",
    x"7B57",
    x"77EE",
    x"73A2",
    x"6E78",
    x"687D",
    x"61BA",
    x"5A3D",
    x"5214",
    x"494F",
    x"3FFE",
    x"3633",
    x"2C01",
    x"217B",
    x"16B5",
    x"0BC4",
    x"00BD",
    x"F5B4",
    x"EABF",
    x"DFF2",
    x"D562",
    x"CB24",
    x"C14A",
    x"B7E8",
    x"AF0F",
    x"A6D0",
    x"9F3C",
    x"985F",
    x"9248",
    x"8D02",
    x"8898",
    x"8510",
    x"8273",
    x"80C5",
    x"800A",
    x"8042",
    x"816E",
    x"838B",
    x"8695",
    x"8A86",
    x"8F57",
    x"94FF",
    x"9B73",
    x"A2A6",
    x"AA8B",
    x"B313",
    x"BC2E",
    x"C5C9",
    x"CFD4",
    x"DA3B",
    x"E4E9",
    x"EFCB",
    x"FACC",
    x"05D7",
    x"10D6",
    x"1BB6",
    x"2661",
    x"30C2",
    x"3AC7",
    x"445C",
    x"4D6F",
    x"55EE",
    x"5DC9",
    x"64F1",
    x"6B5A",
    x"70F6",
    x"75BA",
    x"799E",
    x"7C9B",
    x"7EAA",
    x"7FC8",
    x"7FF2",
    x"7F29",
    x"7D6D",
    x"7AC2",
    x"772E",
    x"72B6",
    x"6D64",
    x"6741",
    x"605A",
    x"58BB",
    x"5073",
    x"4791",
    x"3E28",
    x"3448",
    x"2A04",
    x"1F70",
    x"14A1",
    x"09AA",
    x"FEA1",
    x"F39A",
    x"E8AB",
    x"DDE8",
    x"D366",
    x"C93A",
    x"BF75",
    x"B62C",
    x"AD6F",
    x"A550",
    x"9DDD",
    x"9726",
    x"9136",
    x"8C19",
    x"87D9",
    x"847E",
    x"820E",
    x"808F",
    x"8002",
    x"8069",
    x"81C3",
    x"840D",
    x"8744",
    x"8B61",
    x"905C",
    x"962B",
    x"9CC5",
    x"A41B",
    x"AC20",
    x"B4C6",
    x"BDFA",
    x"C7AD",
    x"D1CA",
    x"DC40",
    x"E6FA",
    x"F1E3",
    x"FCE8",
    x"07F2",
    x"12ED",
    x"1DC4",
    x"2863",
    x"32B4",
    x"3CA5",
    x"4622",
    x"4F1A",
    x"577B",
    x"5F35",
    x"663A",
    x"6C7C",
    x"71F0",
    x"768A",
    x"7A42",
    x"7D12",
    x"7EF3",
    x"7FE3",
    x"7FDE",
    x"7EE6",
    x"7CFD",
    x"7A25",
    x"7664",
    x"71C2",
    x"6C47",
    x"65FE",
    x"5EF3",
    x"5732",
    x"4ECC",
    x"45CF",
    x"3C4D",
    x"3259",
    x"2804",
    x"1D64",
    x"128B",
    x"078F",
    x"FC84",
    x"F180",
    x"E698",
    x"DBE0",
    x"D16E",
    x"C753",
    x"BDA5",
    x"B475",
    x"ABD5",
    x"A3D6",
    x"9C86",
    x"95F3",
    x"902B",
    x"8B38",
    x"8723",
    x"83F5",
    x"81B2",
    x"8061",
    x"8003",
    x"8098",
    x"8220",
    x"8498",
    x"87FC",
    x"8C43",
    x"9168",
    x"975F",
    x"9E1D",
    x"A596",
    x"ADBC",
    x"B67D",
    x"BFCB",
    x"C994",
    x"D3C4",
    x"DE48",
    x"E90D",
    x"F3FD",
    x"FF04",
    x"0A0D",
    x"1503",
    x"1FD1",
    x"2A62",
    x"34A3",
    x"3E7F",
    x"47E4",
    x"50C0",
    x"5902",
    x"609B",
    x"677C",
    x"6D97",
    x"72E2",
    x"7752",
    x"7ADE",
    x"7D81",
    x"7F34",
    x"7FF5",
    x"7FC2",
    x"7E9B",
    x"7C84",
    x"797F",
    x"7593",
    x"70C7",
    x"6B23",
    x"64B4",
    x"5D85",
    x"55A4",
    x"4D1F",
    x"4408",
    x"3A6F",
    x"3066",
    x"2602",
    x"1B55",
    x"1074",
    x"0573",
    x"FA68",
    x"EF68",
    x"E488",
    x"D9DB",
    x"CF78",
    x"C571",
    x"BBD9",
    x"B2C4",
    x"AA41",
    x"A262",
    x"9B35",
    x"94C9",
    x"8F28",
    x"8A5F",
    x"8675",
    x"8374",
    x"815F",
    x"803C",
    x"800C",
    x"80D0",
    x"8287",
    x"852C",
    x"88BC",
    x"8D2E",
    x"927C",
    x"989A",
    x"9F7D",
    x"A718",
    x"AF5C",
    x"B83A",
    x"C1A1",
    x"CB7F",
    x"D5C0",
    x"E053",
    x"EB21",
    x"F617",
    x"0120",
    x"0C27",
    x"1717",
    x"21DB",
    x"2C5F",
    x"368D",
    x"4054",
    x"49A0",
    x"5261",
    x"5A84",
    x"61FA",
    x"68B6",
    x"6EAB",
    x"73CC",
    x"7811",
    x"7B71",
    x"7DE6",
    x"7F6B",
    x"7FFE",
    x"7F9C",
    x"7E48",
    x"7C02",
    x"78D1",
    x"74B9",
    x"6FC3",
    x"69F8",
    x"6363",
    x"5C11",
    x"540F",
    x"4B6D",
    x"423C",
    x"388C",
    x"2E70",
    x"23FC",
    x"1944",
    x"0E5B",
    x"0357",
    x"F84D",
    x"ED51",
    x"E279",
    x"D7D9",
    x"CD86",
    x"C392",
    x"BA12",
    x"B117",
    x"A8B3",
    x"A0F5",
    x"99EC",
    x"93A5",
    x"8E2D",
    x"898E",
    x"85D0",
    x"82FB",
    x"8115",
    x"8020",
    x"801F",
    x"8111",
    x"82F6",
    x"85C8",
    x"8984",
    x"8E21",
    x"9397",
    x"99DC",
    x"A0E3",
    x"A8A0",
    x"B103",
    x"B9FC",
    x"C37B",
    x"CD6D",
    x"D7C0",
    x"E25F",
    x"ED37",
    x"F832",
    x"033D",
    x"0E41",
    x"192A",
    x"23E3",
    x"2E58",
    x"3874",
    x"4225",
    x"4B58",
    x"53FB",
    x"5BFE",
    x"6352",
    x"69E9",
    x"6FB6",
    x"74AE",
    x"78C8",
    x"7BFC",
    x"7E43",
    x"7F9A",
    x"7FFE",
    x"7F6E",
    x"7DEB",
    x"7B78",
    x"781A",
    x"73D7",
    x"6EB8",
    x"68C5",
    x"620B",
    x"5A96",
    x"5275",
    x"49B6",
    x"406B",
    x"36A5",
    x"2C77",
    x"21F5",
    x"1731",
    x"0C42",
    x"013B",
    x"F632",
    x"EB3B",
    x"E06C",
    x"D5D9",
    x"CB97",
    x"C1B8",
    x"B850",
    x"AF71",
    x"A72B",
    x"9F8E",
    x"98A9",
    x"9289",
    x"8D3A",
    x"88C5",
    x"8534",
    x"828C",
    x"80D3",
    x"800D",
    x"803A",
    x"815B",
    x"836E",
    x"866D",
    x"8A54",
    x"8F1C",
    x"94BA",
    x"9B25",
    x"A250",
    x"AA2E",
    x"B2AF",
    x"BBC3",
    x"C559",
    x"CF5F",
    x"D9C2",
    x"E46E",
    x"EF4E",
    x"FA4E",
    x"0559",
    x"1059",
    x"1B3B",
    x"25E8",
    x"304E",
    x"3A57",
    x"43F1",
    x"4D0A",
    x"5590",
    x"5D73",
    x"64A4",
    x"6B15",
    x"70BA",
    x"7588",
    x"7977",
    x"7C7E",
    x"7E98",
    x"7FC0",
    x"7FF5",
    x"7F37",
    x"7D86",
    x"7AE6",
    x"775B",
    x"72EE",
    x"6DA5",
    x"678B",
    x"60AC",
    x"5915",
    x"50D5",
    x"47FA",
    x"3E96",
    x"34BB",
    x"2A7B",
    x"1FEA",
    x"151D",
    x"0A27",
    x"FF1E",
    x"F417",
    x"E927",
    x"DE62",
    x"D3DD",
    x"C9AC",
    x"BFE2",
    x"B693",
    x"ADD0",
    x"A5A9",
    x"9E2E",
    x"976E",
    x"9175",
    x"8C4F",
    x"8805",
    x"849F",
    x"8225",
    x"809B",
    x"8003",
    x"805F",
    x"81AE",
    x"83EE",
    x"871A",
    x"8B2D",
    x"901E",
    x"95E5",
    x"9C75",
    x"A3C4",
    x"ABC1",
    x"B460",
    x"BD8F",
    x"C73C",
    x"D155",
    x"DBC7",
    x"E67E",
    x"F166",
    x"FC6A",
    x"0774",
    x"1271",
    x"1D4A",
    x"27EB",
    -- nota 05
    x"0000",
    x"0BB0",
    x"1746",
    x"22AB",
    x"2DC6",
    x"387F",
    x"42BF",
    x"4C70",
    x"557E",
    x"5DD5",
    x"6564",
    x"6C19",
    x"71E8",
    x"76C2",
    x"7A9F",
    x"7D76",
    x"7F40",
    x"7FFB",
    x"7FA3",
    x"7E3B",
    x"7BC4",
    x"7845",
    x"73C5",
    x"6E4E",
    x"67EA",
    x"60A8",
    x"5898",
    x"4FCA",
    x"4651",
    x"3C42",
    x"31B2",
    x"26B8",
    x"1B6B",
    x"0FE4",
    x"043A",
    x"F888",
    x"ECE5",
    x"E16B",
    x"D633",
    x"CB54",
    x"C0E6",
    x"B6FE",
    x"ADB3",
    x"A518",
    x"9D3F",
    x"9639",
    x"9016",
    x"8AE2",
    x"86A8",
    x"8372",
    x"8146",
    x"8029",
    x"801E",
    x"8124",
    x"8339",
    x"8659",
    x"8A7D",
    x"8F9D",
    x"95AD",
    x"9CA0",
    x"A468",
    x"ACF3",
    x"B631",
    x"C00C",
    x"CA6F",
    x"D546",
    x"E077",
    x"EBED",
    x"F78D",
    x"033F",
    x"0EEA",
    x"1A75",
    x"25C8",
    x"30CA",
    x"3B64",
    x"457E",
    x"4F04",
    x"57E1",
    x"6003",
    x"6756",
    x"6DCD",
    x"7359",
    x"77EF",
    x"7B83",
    x"7E10",
    x"7F8F",
    x"7FFE",
    x"7F5A",
    x"7DA7",
    x"7AE6",
    x"771F",
    x"7259",
    x"6C9F",
    x"65FC",
    x"5E7F",
    x"5639",
    x"4D39",
    x"4395",
    x"3960",
    x"2EB0",
    x"239D",
    x"183D",
    x"0CAA",
    x"00FB",
    x"F54B",
    x"E9B1",
    x"DE47",
    x"D325",
    x"C863",
    x"BE18",
    x"B45A",
    x"AB3E",
    x"A2D7",
    x"9B37",
    x"946E",
    x"8E8C",
    x"899C",
    x"85AA",
    x"82BD",
    x"80DC",
    x"800B",
    x"804B",
    x"819D",
    x"83FC",
    x"8765",
    x"8BD0",
    x"9134",
    x"9784",
    x"9EB4",
    x"A6B4",
    x"AF72",
    x"B8DD",
    x"C2E1",
    x"CD66",
    x"D858",
    x"E39F",
    x"EF23",
    x"FACB",
    x"067D",
    x"1222",
    x"1DA0",
    x"28DF",
    x"33C6",
    x"3E3F",
    x"4832",
    x"518C",
    x"5A36",
    x"6220",
    x"6938",
    x"6F6F",
    x"74B8",
    x"7907",
    x"7C53",
    x"7E96",
    x"7FC9",
    x"7FEC",
    x"7EFD",
    x"7CFE",
    x"79F4",
    x"75E5",
    x"70DB",
    x"6ADE",
    x"63FE",
    x"5C47",
    x"53CB",
    x"4A9C",
    x"40CE",
    x"3675",
    x"2BA7",
    x"207C",
    x"150C",
    x"096E",
    x"FDBC",
    x"F210",
    x"E681",
    x"DB28",
    x"D01F",
    x"C57B",
    x"BB55",
    x"B1C2",
    x"A8D6",
    x"A0A4",
    x"993F",
    x"92B5",
    x"8D15",
    x"886A",
    x"84BF",
    x"821C",
    x"8086",
    x"8001",
    x"808D",
    x"822A",
    x"84D4",
    x"8886",
    x"8D37",
    x"92DD",
    x"996D",
    x"A0D8",
    x"A90E",
    x"B1FF",
    x"BB96",
    x"C5C0",
    x"D066",
    x"DB72",
    x"E6CC",
    x"F25C",
    x"FE09",
    x"09BB",
    x"1557",
    x"20C6",
    x"2BEF",
    x"36BA",
    x"4110",
    x"4ADB",
    x"5405",
    x"5C7C",
    x"642E",
    x"6B09",
    x"70FF",
    x"7603",
    x"7A0B",
    x"7D0F",
    x"7F06",
    x"7FEE",
    x"7FC5",
    x"7E8A",
    x"7C41",
    x"78EE",
    x"7498",
    x"6F49",
    x"690C",
    x"61EF",
    x"5A00",
    x"5150",
    x"47F3",
    x"3DFC",
    x"3380",
    x"2896",
    x"1D56",
    x"11D6",
    x"0631",
    x"FA7E",
    x"EED7",
    x"E355",
    x"D810",
    x"CD20",
    x"C29D",
    x"B89E",
    x"AF37",
    x"A67D",
    x"9E82",
    x"9758",
    x"910D",
    x"8BB0",
    x"874C",
    x"83EA",
    x"8191",
    x"8046",
    x"800D",
    x"80E5",
    x"82CD",
    x"85C0",
    x"89BA",
    x"8EB0",
    x"9498",
    x"9B66",
    x"A30B",
    x"AB77",
    x"B498",
    x"BE5A",
    x"C8A8",
    x"D36D",
    x"DE91",
    x"E9FD",
    x"F597",
    x"0148",
    x"0CF6",
    x"1889",
    x"23E7",
    x"2EF8",
    x"39A5",
    x"43D6",
    x"4D76",
    x"5671",
    x"5EB3",
    x"662B",
    x"6CC7",
    x"727C",
    x"773B",
    x"7AFC",
    x"7DB5",
    x"7F62",
    x"7FFE",
    x"7F89",
    x"7E03",
    x"7B6F",
    x"77D4",
    x"7338",
    x"6DA6",
    x"6729",
    x"5FD0",
    x"57AA",
    x"4EC8",
    x"453E",
    x"3B20",
    x"3083",
    x"257F",
    x"1A2A",
    x"0E9E",
    x"02F2",
    x"F740",
    x"EBA1",
    x"E02D",
    x"D4FD",
    x"CA2A",
    x"BFC9",
    x"B5F2",
    x"ACB9",
    x"A432",
    x"9C70",
    x"9582",
    x"8F78",
    x"8A5F",
    x"8641",
    x"8328",
    x"811A",
    x"801B",
    x"802D",
    x"8151",
    x"8384",
    x"86C1",
    x"8B01",
    x"903B",
    x"9665",
    x"9D70",
    x"A54E",
    x"ADEE",
    x"B73E",
    x"C129",
    x"CB9A",
    x"D67C",
    x"E1B6",
    x"ED31",
    x"F8D4",
    x"0487",
    x"1030",
    x"1BB6",
    x"2701",
    x"31F9",
    x"3C86",
    x"4691",
    x"5006",
    x"58CF",
    x"60DA",
    x"6817",
    x"6E74",
    x"73E6",
    x"7860",
    x"7BD8",
    x"7E47",
    x"7FA9",
    x"7FF9",
    x"7F38",
    x"7D67",
    x"7A89",
    x"76A6",
    x"71C4",
    x"6BF0",
    x"6535",
    x"5DA1",
    x"5545",
    x"4C33",
    x"427D",
    x"383A",
    x"2D7E",
    x"2261",
    x"16FB",
    x"0B63",
    x"FFB3",
    x"F404",
    x"E86E",
    x"DD0B",
    x"D1F2",
    x"C73C",
    x"BD00",
    x"B352",
    x"AA49",
    x"A1F7",
    x"9A6E",
    x"93BE",
    x"8DF6",
    x"8921",
    x"854B",
    x"827B",
    x"80B8",
    x"8004",
    x"8063",
    x"81D2",
    x"844F",
    x"87D5",
    x"8C5C",
    x"91D9",
    x"9843",
    x"9F8A",
    x"A7A0",
    x"B072",
    x"B9EF",
    x"C402",
    x"CE94",
    x"D991",
    x"E4E0",
    x"F068",
    x"FC12",
    x"07C5",
    x"1367",
    x"1EDF",
    x"2A15",
    x"34F2",
    x"3F5D",
    x"4940",
    x"5287",
    x"5B1E",
    x"62F2",
    x"69F2",
    x"700F",
    x"753D",
    x"7970",
    x"7CA0",
    x"7EC5",
    x"7FDA",
    x"7FDF",
    x"7ED2",
    x"7CB6",
    x"798F",
    x"7564",
    x"703E",
    x"6A29",
    x"6330",
    x"5B63",
    x"52D2",
    x"4991",
    x"3FB2",
    x"354B",
    x"2A72",
    x"1F3E",
    x"13C8",
    x"0827",
    x"FC74",
    x"F0CA",
    x"E540",
    x"D9EF",
    x"CEEF",
    x"C458",
    x"BA41",
    x"B0BF",
    x"A7E7",
    x"9FCB",
    x"987C",
    x"920C",
    x"8C86",
    x"87F7",
    x"8469",
    x"81E3",
    x"806A",
    x"8003",
    x"80AD",
    x"8268",
    x"852F",
    x"88FD",
    x"8DC9",
    x"938A",
    x"9A32",
    x"A1B4",
    x"AA00",
    x"B304",
    x"BCAC",
    x"C6E5",
    x"D197",
    x"DCAD",
    x"E80E",
    x"F3A2",
    x"FF51",
    x"0B02",
    x"169A",
    x"2203",
    x"2D23",
    x"37E2",
    x"422A",
    x"4BE4",
    x"54FC",
    x"5D5E",
    x"64F9",
    x"6BBB",
    x"7197",
    x"7681",
    x"7A6D",
    x"7D53",
    x"7F2D",
    x"7FF7",
    x"7FB0",
    x"7E57",
    x"7BF1",
    x"7881",
    x"740F",
    x"6EA6",
    x"6850",
    x"611A",
    x"5915",
    x"5052",
    x"46E3",
    x"3CDC",
    x"3253",
    x"275F",
    x"1C16",
    x"1091",
    x"04E9",
    x"F936",
    x"ED92",
    x"E215",
    x"D6D8",
    x"CBF4",
    x"C17E",
    x"B78E",
    x"AE39",
    x"A593",
    x"9DAF",
    x"969C",
    x"906B",
    x"8B29",
    x"86E0",
    x"839B",
    x"815F",
    x"8032",
    x"8017",
    x"810D",
    x"8312",
    x"8623",
    x"8A38",
    x"8F4A",
    x"954C",
    x"9C32",
    x"A3EE",
    x"AC6F",
    x"B5A2",
    x"BF74",
    x"C9D1",
    x"D4A1",
    x"DFCE",
    x"EB40",
    x"F6DE",
    x"0290",
    x"0E3D",
    x"19CA",
    x"2521",
    x"3028",
    x"3AC9",
    x"44EB",
    x"4E7B",
    x"5762",
    x"5F8F",
    x"66EF",
    x"6D73",
    x"730D",
    x"77B1",
    x"7B55",
    x"7DF1",
    x"7F80",
    x"7FFF",
    x"7F6B",
    x"7DC8",
    x"7B17",
    x"775F",
    x"72A7",
    x"6CFB",
    x"6665",
    x"5EF5",
    x"56B9",
    x"4DC4",
    x"4429",
    x"39FC",
    x"2F53",
    x"2445",
    x"18E9",
    x"0D58",
    x"01AA",
    x"F5F9",
    x"EA5D",
    x"DEF0",
    x"D3C9",
    x"C901",
    x"BEAE",
    x"B4E7",
    x"ABC1",
    x"A34F",
    x"9BA3",
    x"94CD",
    x"8EDD",
    x"89DF",
    x"85DE",
    x"82E1",
    x"80F0",
    x"800F",
    x"8040",
    x"8181",
    x"83D2",
    x"872B",
    x"8B87",
    x"90DD",
    x"971F",
    x"9E43",
    x"A637",
    x"AEEB",
    x"B84C",
    x"C247",
    x"CCC6",
    x"D7B3",
    x"E2F5",
    x"EE76",
    x"FA1C",
    x"05CF",
    x"1175",
    x"1CF6",
    x"2839",
    x"3326",
    x"3DA6",
    x"47A2",
    x"5105",
    x"59BA",
    x"61B0",
    x"68D4",
    x"6F19",
    x"7470",
    x"78CE",
    x"7C29",
    x"7E7B",
    x"7FBF",
    x"7FF1",
    x"7F12",
    x"7D23",
    x"7A29",
    x"7629",
    x"712D",
    x"6B3E",
    x"646A",
    x"5CC0",
    x"544F",
    x"4B2A",
    x"4164",
    x"3713",
    x"2C4B",
    x"2125",
    x"15B8",
    x"0A1C",
    x"FE6B",
    x"F2BD",
    x"E72C",
    x"DBD0",
    x"D0C1",
    x"C617",
    x"BBE9",
    x"B24D",
    x"A956",
    x"A119",
    x"99A7",
    x"9310",
    x"8D62",
    x"88A9",
    x"84EF",
    x"823C",
    x"8097",
    x"8001",
    x"807E",
    x"820B",
    x"84A5",
    x"8847",
    x"8CEA",
    x"9282",
    x"9904",
    x"A063",
    x"A88E",
    x"B174",
    x"BB03",
    x"C524",
    x"CFC4",
    x"DACA",
    x"E621",
    x"F1AE",
    x"FD5A",
    x"090C",
    x"14AB",
    x"201D",
    x"2B4B",
    x"361C",
    x"4079",
    x"4A4D",
    x"5381",
    x"5C03",
    x"63C0",
    x"6AA8",
    x"70AC",
    x"75BF",
    x"79D6",
    x"7CE9",
    x"7EF0",
    x"7FE8",
    x"7FCF",
    x"7EA4",
    x"7C6A",
    x"7927",
    x"74E0",
    x"6F9F",
    x"6970",
    x"625F",
    x"5A7C",
    x"51D7",
    x"4883",
    x"3E95",
    x"3420",
    x"293C",
    x"1E00",
    x"1283",
    x"06DF",
    x"FB2C",
    x"EF84",
    x"E3FF",
    x"D8B6",
    x"CDC1",
    x"C337",
    x"B92F",
    x"AFBF",
    x"A6FA",
    x"9EF4",
    x"97BD",
    x"9165",
    x"8BFA",
    x"8786",
    x"8415",
    x"81AC",
    x"8052",
    x"8008",
    x"80D1",
    x"82A9",
    x"858D",
    x"8977",
    x"8E5F",
    x"9439",
    x"9AFA",
    x"A293",
    x"AAF4",
    x"B40B",
    x"BDC4",
    x"C80B",
    x"D2C9",
    x"DDE9",
    x"E951",
    x"F4E9",
    x"0099",
    x"0C48",
    x"17DD",
    x"233F",
    x"2E55",
    x"3908",
    x"4342",
    x"4CEB",
    x"55F0",
    x"5E3D",
    x"65C1",
    x"6C6B",
    x"722D",
    x"76FB",
    x"7ACB",
    x"7D94",
    x"7F50",
    x"7FFD",
    x"7F97",
    x"7E21",
    x"7B9D",
    x"7811",
    x"7384",
    x"6DFF",
    x"6790",
    x"6043",
    x"5829",
    x"4F51",
    x"45D1",
    x"3BBB",
    x"3125",
    x"2626",
    x"1AD5",
    x"0F4B",
    x"03A1",
    x"F7EF",
    x"EC4E",
    x"E0D7",
    x"D5A2",
    x"CAC8",
    x"C061",
    x"B681",
    x"AD3E",
    x"A4AC",
    x"9CDE",
    x"95E3",
    x"8FCC",
    x"8AA4",
    x"8678",
    x"834F",
    x"8131",
    x"8022",
    x"8025",
    x"8138",
    x"835C",
    x"8689",
    x"8ABA",
    x"8FE7",
    x"9602",
    x"9D01",
    x"A4D3",
    x"AD68",
    x"B6AE",
    x"C091",
    x"CAFB",
    x"D5D6",
    x"E10C",
    x"EC84",
    x"F826",
    x"03D8",
    x"0F82",
    x"1B0B",
    x"265B",
    x"3158",
    x"3BEB",
    x"45FF",
    x"4F7D",
    x"5851",
    x"6068",
    x"67B1",
    x"6E1C",
    x"739B",
    x"7824",
    x"7BAB",
    x"7E2A",
    x"7F9C",
    x"7FFC",
    x"7F4B",
    x"7D89",
    x"7ABB",
    x"76E7",
    x"7214",
    x"6C4E",
    x"659F",
    x"5E18",
    x"55C7",
    x"4CBF",
    x"4312",
    x"38D7",
    x"2E21",
    x"230A",
    x"17A7",
    x"0C11",
    x"0062",
    x"F4B2",
    x"E91A",
    x"DDB3",
    x"D296",
    x"C7D9",
    x"BD95",
    x"B3DE",
    x"AACB",
    x"A26E",
    x"9AD8",
    x"941C",
    x"8E45",
    x"8962",
    x"857D",
    x"829E",
    x"80CA",
    x"8007",
    x"8056",
    x"81B5",
    x"8423",
    x"8799",
    x"8C11",
    x"9181",
    x"97DD",
    x"9F18",
    x"A722",
    x"AFEA",
    x"B95D",
    x"C368",
    x"CDF3",
    x"D8EA",
    x"E435",
    x"EFBB",
    x"FB64",
    x"0716",
    x"12BA",
    x"1E35",
    x"2970",
    x"3452",
    x"3EC5",
    x"48B1",
    x"5202",
    x"5AA3",
    x"6282",
    x"698F",
    x"6FBA",
    x"74F6",
    x"7938",
    x"7C77",
    x"7EAC",
    x"7FD2",
    x"7FE6",
    x"7EE9",
    x"7CDD",
    x"79C5",
    x"75A9",
    x"7092",
    x"6A8A",
    x"639E",
    x"5BDD",
    x"5357",
    x"4A20",
    x"4049",
    x"35EA",
    x"2B17",
    x"1FE8",
    x"1474",
    x"08D5",
    x"FD23",
    x"F177",
    x"E5EB",
    x"DA96",
    x"CF91",
    x"C4F3",
    x"BAD4",
    x"B149",
    x"A866",
    x"A03E",
    x"98E4",
    x"9265",
    x"8CD1",
    x"8834",
    x"8496",
    x"8201",
    x"8079",
    x"8002",
    x"809C",
    x"8247",
    x"84FE",
    x"88BD",
    x"8D7B",
    x"932D",
    x"99C9",
    x"A13F",
    x"A97F",
    x"B279",
    x"BC18",
    x"C648",
    x"D0F4",
    x"DC05",
    x"E762",
    x"F2F4",
    x"FEA3",
    x"0A53",
    x"15EE",
    x"215A",
    x"2C7F",
    x"3744",
    x"4194",
    x"4B57",
    x"5479",
    x"5CE6",
    x"648D",
    x"6B5C",
    x"7146",
    x"763E",
    x"7A39",
    x"7D2F",
    x"7F19",
    x"7FF3",
    x"7FBB",
    x"7E73",
    x"7C1C",
    x"78BB",
    x"7459",
    x"6EFD",
    x"68B4",
    x"618C",
    x"5993",
    x"50DA",
    x"4774",
    x"3D76",
    x"32F4",
    x"2805",
    x"1CC0",
    x"113E",
    x"0597",
    x"F9E5",
    x"EE3F",
    x"E2BF",
    x"D77E",
    x"CC93",
    x"C217",
    x"B81F",
    x"AEC0",
    x"A60F",
    x"9E1F",
    x"9700",
    x"90C1",
    x"8B71",
    x"8719",
    x"83C4",
    x"8179",
    x"803C",
    x"8011",
    x"80F7",
    x"82ED",
    x"85EE",
    x"89F4",
    x"8EF7",
    x"94EC",
    x"9BC5",
    x"A375",
    x"ABEB",
    -- nota 06
    x"0000",
    x"0C61",
    x"18A4",
    x"24AC",
    x"305C",
    x"3B98",
    x"4645",
    x"504A",
    x"598D",
    x"61FA",
    x"697C",
    x"7000",
    x"7578",
    x"79D5",
    x"7D0F",
    x"7F1C",
    x"7FF8",
    x"7FA1",
    x"7E17",
    x"7B5F",
    x"777F",
    x"7280",
    x"6C6F",
    x"6559",
    x"5D50",
    x"5466",
    x"4AB3",
    x"404C",
    x"354A",
    x"29C9",
    x"1DE4",
    x"11B7",
    x"055F",
    x"F8FA",
    x"ECA7",
    x"E081",
    x"D4A7",
    x"C936",
    x"BE48",
    x"B3F7",
    x"AA5D",
    x"A191",
    x"99A7",
    x"92B3",
    x"8CC5",
    x"87EC",
    x"8433",
    x"81A3",
    x"8042",
    x"8014",
    x"8119",
    x"834E",
    x"86AF",
    x"8B33",
    x"90CF",
    x"9776",
    x"9F18",
    x"A7A3",
    x"B102",
    x"BB1E",
    x"C5E0",
    x"D12D",
    x"DCEA",
    x"E8FC",
    x"F545",
    x"01A7",
    x"0E06",
    x"1A43",
    x"2641",
    x"31E3",
    x"3D0E",
    x"47A6",
    x"5192",
    x"5ABA",
    x"6308",
    x"6A69",
    x"70CB",
    x"761D",
    x"7A55",
    x"7D66",
    x"7F4B",
    x"7FFE",
    x"7F7E",
    x"7DCC",
    x"7AEC",
    x"76E5",
    x"71C1",
    x"6B8B",
    x"6454",
    x"5C2C",
    x"5326",
    x"4959",
    x"3EDC",
    x"33C8",
    x"2838",
    x"1C48",
    x"1013",
    x"03B8",
    x"F754",
    x"EB04",
    x"DEE8",
    x"D31A",
    x"C7B8",
    x"BCDE",
    x"B2A4",
    x"A924",
    x"A075",
    x"98AB",
    x"91D9",
    x"8C0F",
    x"875C",
    x"83CA",
    x"8162",
    x"802A",
    x"8025",
    x"8153",
    x"83B0",
    x"8739",
    x"8BE3",
    x"91A3",
    x"986D",
    x"A02F",
    x"A8D7",
    x"B250",
    x"BC84",
    x"C75A",
    x"D2B8",
    x"DE82",
    x"EA9D",
    x"F6EB",
    x"034F",
    x"0FAB",
    x"1BE1",
    x"27D4",
    x"3368",
    x"3E81",
    x"4903",
    x"52D6",
    x"5BE3",
    x"6412",
    x"6B52",
    x"7190",
    x"76BE",
    x"7ACE",
    x"7DB8",
    x"7F74",
    x"7FFF",
    x"7F56",
    x"7D7B",
    x"7A73",
    x"7646",
    x"70FC",
    x"6AA4",
    x"634B",
    x"5B04",
    x"51E3",
    x"47FD",
    x"3D6A",
    x"3244",
    x"26A5",
    x"1AAA",
    x"0E6F",
    x"0211",
    x"F5AE",
    x"E963",
    x"DD4F",
    x"D18F",
    x"C63D",
    x"BB77",
    x"B155",
    x"A7EF",
    x"9F5D",
    x"97B3",
    x"9104",
    x"8B5E",
    x"86D1",
    x"8366",
    x"8127",
    x"8018",
    x"803B",
    x"8192",
    x"8418",
    x"87C7",
    x"8C97",
    x"927C",
    x"9968",
    x"A14A",
    x"AA0F",
    x"B3A3",
    x"BDED",
    x"C8D7",
    x"D445",
    x"E01B",
    x"EC3E",
    x"F891",
    x"04F6",
    x"114E",
    x"1D7D",
    x"2966",
    x"34EB",
    x"3FF1",
    x"4A5D",
    x"5417",
    x"5D07",
    x"6518",
    x"6C37",
    x"7251",
    x"7759",
    x"7B43",
    x"7E05",
    x"7F99",
    x"7FFA",
    x"7F28",
    x"7D25",
    x"79F5",
    x"75A1",
    x"7033",
    x"69B7",
    x"623E",
    x"59D8",
    x"509C",
    x"469D",
    x"3BF5",
    x"30BE",
    x"2511",
    x"190B",
    x"0CCA",
    x"0069",
    x"F408",
    x"E7C3",
    x"DBB9",
    x"D005",
    x"C4C5",
    x"BA13",
    x"B008",
    x"A6BE",
    x"9E4A",
    x"96C0",
    x"9033",
    x"8AB2",
    x"864B",
    x"8308",
    x"80F1",
    x"800B",
    x"8057",
    x"81D7",
    x"8485",
    x"885B",
    x"8D51",
    x"935A",
    x"9A67",
    x"A269",
    x"AB4B",
    x"B4F8",
    x"BF59",
    x"CA56",
    x"D5D3",
    x"E1B6",
    x"EDE1",
    x"FA38",
    x"069D",
    x"12F1",
    x"1F19",
    x"2AF5",
    x"366B",
    x"415E",
    x"4BB4",
    x"5555",
    x"5E28",
    x"661A",
    x"6D16",
    x"730D",
    x"77F0",
    x"7BB3",
    x"7E4C",
    x"7FB7",
    x"7FF0",
    x"7EF5",
    x"7CC9",
    x"7972",
    x"74F8",
    x"6F65",
    x"68C6",
    x"612C",
    x"58A9",
    x"4F51",
    x"453B",
    x"3A7E",
    x"2F35",
    x"237B",
    x"176C",
    x"0B24",
    x"FEC2",
    x"F263",
    x"E624",
    x"DA23",
    x"CE7E",
    x"C34F",
    x"B8B2",
    x"AEC0",
    x"A590",
    x"9D3A",
    x"95D1",
    x"8F67",
    x"8A0B",
    x"85CB",
    x"82AF",
    x"80C0",
    x"8003",
    x"8079",
    x"8221",
    x"84F7",
    x"88F4",
    x"8E0F",
    x"943C",
    x"9B6B",
    x"A38B",
    x"AC8A",
    x"B650",
    x"C0C8",
    x"CBD7",
    x"D764",
    x"E352",
    x"EF85",
    x"FBDF",
    x"0843",
    x"1494",
    x"20B3",
    x"2C83",
    x"37E9",
    x"42C9",
    x"4D08",
    x"568E",
    x"5F45",
    x"6717",
    x"6DF1",
    x"73C4",
    x"7881",
    x"7C1D",
    x"7E8F",
    x"7FD1",
    x"7FE0",
    x"7EBC",
    x"7C68",
    x"78EA",
    x"744A",
    x"6E92",
    x"67D1",
    x"6017",
    x"5776",
    x"4E03",
    x"43D5",
    x"3904",
    x"2DAB",
    x"21E4",
    x"15CB",
    x"097E",
    x"FD1B",
    x"F0BE",
    x"E486",
    x"D890",
    x"CCF8",
    x"C1DB",
    x"B754",
    x"AD7A",
    x"A467",
    x"9C2F",
    x"94E7",
    x"8EA0",
    x"896A",
    x"854F",
    x"825C",
    x"8095",
    x"8001",
    x"80A0",
    x"8270",
    x"856E",
    x"8992",
    x"8ED2",
    x"9522",
    x"9C73",
    x"A4B2",
    x"ADCC",
    x"B7AC",
    x"C23A",
    x"CD5B",
    x"D8F6",
    x"E4EF",
    x"F129",
    x"FD86",
    x"09EA",
    x"1635",
    x"224B",
    x"2E0F",
    x"3965",
    x"4430",
    x"4E58",
    x"57C4",
    x"605E",
    x"6810",
    x"6EC8",
    x"7476",
    x"790D",
    x"7C82",
    x"7ECB",
    x"7FE4",
    x"7FCB",
    x"7E7E",
    x"7C02",
    x"785D",
    x"7396",
    x"6DBA",
    x"66D7",
    x"5EFD",
    x"563F",
    x"4CB2",
    x"426D",
    x"3788",
    x"2C1E",
    x"204B",
    x"1429",
    x"07D8",
    x"FB73",
    x"EF1A",
    x"E2E9",
    x"D6FE",
    x"CB75",
    x"C06B",
    x"B5F9",
    x"AC38",
    x"A341",
    x"9B28",
    x"9402",
    x"8DDE",
    x"88CD",
    x"84D9",
    x"820E",
    x"8070",
    x"8004",
    x"80CC",
    x"82C5",
    x"85EB",
    x"8A35",
    x"8F9B",
    x"960E",
    x"9D7F",
    x"A5DD",
    x"AF13",
    x"B90B",
    x"C3AE",
    x"CEE1",
    x"DA8A",
    x"E68D",
    x"F2CE",
    x"FF2D",
    x"0B8F",
    x"17D5",
    x"23E2",
    x"2F99",
    x"3ADE",
    x"4595",
    x"4FA5",
    x"58F6",
    x"6172",
    x"6904",
    x"6F9A",
    x"7523",
    x"7994",
    x"7CE1",
    x"7F02",
    x"7FF3",
    x"7FB0",
    x"7E3B",
    x"7B97",
    x"77CA",
    x"72DE",
    x"6CDE",
    x"65D9",
    x"5DDF",
    x"5504",
    x"4B5D",
    x"4101",
    x"360A",
    x"2A90",
    x"1EB0",
    x"1287",
    x"0631",
    x"F9CD",
    x"ED77",
    x"E14D",
    x"D56E",
    x"C9F4",
    x"BEFD",
    x"B4A1",
    x"AAFA",
    x"A21F",
    x"9A26",
    x"9321",
    x"8D21",
    x"8835",
    x"8469",
    x"81C5",
    x"8050",
    x"800D",
    x"80FE",
    x"831F",
    x"866D",
    x"8ADE",
    x"9068",
    x"96FD",
    x"9E8F",
    x"A70B",
    x"B05C",
    x"BA6D",
    x"C524",
    x"D069",
    x"DC20",
    x"E82D",
    x"F473",
    x"00D5",
    x"0D35",
    x"1975",
    x"2578",
    x"3121",
    x"3C54",
    x"46F7",
    x"50EF",
    x"5A25",
    x"6283",
    x"69F4",
    x"7066",
    x"75CC",
    x"7A16",
    x"7D3B",
    x"7F34",
    x"7FFC",
    x"7F90",
    x"7DF2",
    x"7B26",
    x"7732",
    x"7221",
    x"6BFD",
    x"64D6",
    x"5CBD",
    x"53C6",
    x"4A05",
    x"3F93",
    x"3489",
    x"2900",
    x"1D15",
    x"10E4",
    x"048A",
    x"F826",
    x"EBD4",
    x"DFB3",
    x"D3DF",
    x"C876",
    x"BD91",
    x"B34C",
    x"A9BF",
    x"A102",
    x"9928",
    x"9245",
    x"8C69",
    x"87A3",
    x"83FD",
    x"8181",
    x"8035",
    x"801C",
    x"8135",
    x"837F",
    x"86F4",
    x"8B8B",
    x"9139",
    x"97F2",
    x"9FA4",
    x"A83D",
    x"B1AA",
    x"BBD2",
    x"C69D",
    x"D1F3",
    x"DDB7",
    x"E9CD",
    x"F619",
    x"027C",
    x"0EDA",
    x"1B13",
    x"270C",
    x"32A7",
    x"3DC9",
    x"4856",
    x"5235",
    x"5B50",
    x"638F",
    x"6ADF",
    x"712F",
    x"766F",
    x"7A92",
    x"7D90",
    x"7F60",
    x"7FFF",
    x"7F6A",
    x"7DA4",
    x"7AB0",
    x"7696",
    x"715F",
    x"6B17",
    x"63CF",
    x"5B98",
    x"5284",
    x"48AB",
    x"3E23",
    x"3306",
    x"276E",
    x"1B78",
    x"0F40",
    x"02E3",
    x"F67F",
    x"EA33",
    x"DE1A",
    x"D253",
    x"C6FA",
    x"BC29",
    x"B1FB",
    x"A888",
    x"9FE8",
    x"982E",
    x"916D",
    x"8BB6",
    x"8715",
    x"8397",
    x"8143",
    x"8020",
    x"8030",
    x"8172",
    x"83E4",
    x"8780",
    x"8C3D",
    x"9210",
    x"98EA",
    x"A0BD",
    x"A973",
    x"B2FA",
    x"BD39",
    x"C819",
    x"D37F",
    x"DF50",
    x"EB6F",
    x"F7BF",
    x"0423",
    x"107E",
    x"1CB0",
    x"289E",
    x"342B",
    x"3F3A",
    x"49B1",
    x"5378",
    x"5C76",
    x"6497",
    x"6BC6",
    x"71F2",
    x"770D",
    x"7B0A",
    x"7DE0",
    x"7F87",
    x"7FFD",
    x"7F3F",
    x"7D50",
    x"7A35",
    x"75F4",
    x"7098",
    x"6A2D",
    x"62C4",
    x"5A6E",
    x"513F",
    x"474C",
    x"3CAF",
    x"3180",
    x"25DA",
    x"19DA",
    x"0D9B",
    x"013C",
    x"F4D9",
    x"E892",
    x"DC83",
    x"D0C9",
    x"C580",
    x"BAC3",
    x"B0AD",
    x"A755",
    x"9ED2",
    x"9738",
    x"909A",
    x"8B07",
    x"868D",
    x"8336",
    x"810B",
    x"8010",
    x"8049",
    x"81B4",
    x"844E",
    x"8811",
    x"8CF4",
    x"92EB",
    x"99E8",
    x"A1D9",
    x"AAAD",
    x"B44E",
    x"BEA4",
    x"C997",
    x"D50D",
    x"E0EA",
    x"ED11",
    x"F966",
    x"05CA",
    x"1221",
    x"1E4C",
    x"2A2F",
    x"35AC",
    x"40A9",
    x"4B0A",
    x"54B7",
    x"5D99",
    x"659A",
    x"6CA8",
    x"72B0",
    x"77A6",
    x"7B7C",
    x"7E2A",
    x"7FA9",
    x"7FF5",
    x"7F0F",
    x"7CF8",
    x"79B4",
    x"754D",
    x"6FCC",
    x"693F",
    x"61B5",
    x"5940",
    x"4FF6",
    x"45EB",
    x"3B39",
    x"2FF9",
    x"2445",
    x"183B",
    x"0BF6",
    x"FF94",
    x"F334",
    x"E6F2",
    x"DAED",
    x"CF40",
    x"C408",
    x"B961",
    x"AF63",
    x"A626",
    x"9DC1",
    x"9648",
    x"8FCC",
    x"8A5E",
    x"860A",
    x"82DB",
    x"80D8",
    x"8006",
    x"8068",
    x"81FB",
    x"84BD",
    x"88A7",
    x"8DB0",
    x"93CB",
    x"9AE9",
    x"A2FA",
    x"ABEB",
    x"B5A5",
    x"C011",
    x"CB17",
    x"D69C",
    x"E285",
    x"EEB4",
    x"FB0D",
    x"0771",
    x"13C4",
    x"1FE7",
    x"2BBE",
    x"372B",
    x"4215",
    x"4C5F",
    x"55F3",
    x"5EB8",
    x"669A",
    x"6D85",
    x"736A",
    x"7839",
    x"7BE9",
    x"7E6E",
    x"7FC5",
    x"7FE8",
    x"7ED9",
    x"7C99",
    x"792E",
    x"74A1",
    x"6EFB",
    x"684B",
    x"60A1",
    x"580F",
    x"4EAA",
    x"4487",
    x"39C1",
    x"2E6F",
    x"22AE",
    x"169A",
    x"0A50",
    x"FDED",
    x"F18F",
    x"E554",
    x"D958",
    x"CDBA",
    x"C294",
    x"B801",
    x"AE1C",
    x"A4FA",
    x"9CB4",
    x"955B",
    x"8F03",
    x"89B9",
    x"858C",
    x"8284",
    x"80AA",
    x"8001",
    x"808C",
    x"8248",
    x"8532",
    x"8943",
    x"8E71",
    x"94AF",
    x"9BEF",
    x"A41F",
    x"AD2C",
    x"B6FF",
    x"C181",
    x"CC9A",
    x"D82E",
    x"E421",
    x"F058",
    x"FCB4",
    x"0918",
    x"1566",
    x"2180",
    x"2D4B",
    x"38A8",
    x"437E",
    x"4DB1",
    x"572B",
    x"5FD2",
    x"6794",
    x"6E5E",
    x"741E",
    x"78C8",
    x"7C50",
    x"7EAE",
    x"7FDB",
    x"7FD6",
    x"7E9E",
    x"7C36",
    x"78A4",
    x"73F0",
    x"6E26",
    x"6754",
    x"5F8A",
    x"56DA",
    x"4D5A",
    x"4320",
    x"3846",
    x"2CE4",
    x"2116",
    x"14F9",
    x"08AA",
    x"FC46",
    x"EFEB",
    x"E3B6",
    x"D7C6",
    x"CC35",
    x"C122",
    x"B6A5",
    x"ACD8",
    x"A3D3",
    x"9BAB",
    x"9473",
    x"8E3E",
    x"891A",
    x"8513",
    x"8234",
    x"8082",
    x"8002",
    x"80B5",
    x"829A",
    x"85AC",
    x"89E4",
    x"8F37",
    x"9598",
    x"9CF9",
    x"A548",
    x"AE70",
    x"B85C",
    x"C2F4",
    x"CE1F",
    x"D9C1",
    x"E5BF",
    x"F1FC",
    x"FE5B",
    x"0ABE",
    x"1707",
    x"2318",
    x"2ED6",
    x"3A23",
    x"44E4",
    x"4F00",
    x"585F",
    x"60E9",
    x"688B",
    x"6F32",
    x"74CE",
    x"7952",
    x"7CB2",
    x"7EE8",
    x"7FEC",
    x"7FBE",
    x"7E5D",
    x"7BCD",
    x"7814",
    x"733A",
    x"6D4C",
    x"6658",
    x"5E6E",
    x"55A1",
    x"4C07",
    x"41B6",
    x"36C8",
    x"2B56",
    x"1F7D",
    x"1357",
    x"0703",
    x"FA9F",
    x"EE47",
    x"E21A",
    x"D635",
    x"CAB3",
    x"BFB2",
    x"B54B",
    x"AB98",
    x"A2AF",
    x"9AA6",
    x"9390",
    x"8D7F",
    x"8880",
    x"84A0",
    x"81E8",
    x"805F",
    x"8008",
    x"80E5",
    x"82F2",
    x"862B",
    x"8A89",
    x"9001",
    x"9686",
    x"9E07",
    x"A674",
    x"AFB8",
    x"B9BD",
    x"C46A",
    x"CFA6",
    x"DB56",
    x"E75E",
    x"F3A1",
    x"0002",
    x"0C63",
    x"18A6",
    x"24AF",
    x"305F",
    x"3B9A",
    x"4647",
    x"504C",
    x"598F",
    x"61FC",
    x"697D",
    x"7001",
    x"7579",
    x"79D6",
    x"7D0F",
    x"7F1C",
    x"7FF8",
    x"7FA1",
    x"7E17",
    x"7B5F",
    x"777E",
    x"727F",
    x"6C6D",
    x"6557",
    x"5D4E",
    x"5465",
    x"4AB1",
    x"404A",
    x"3548",
    x"29C7",
    x"1DE2",
    x"11B4",
    x"055D",
    x"F8F8",
    x"ECA4",
    x"E07F",
    x"D4A5",
    x"C934",
    x"BE46",
    x"B3F5",
    x"AA5B",
    x"A18F",
    x"99A6",
    x"92B2",
    x"8CC4",
    x"87EB",
    x"8432",
    x"81A2",
    x"8042",
    x"8014",
    x"8119",
    -- nota 07
    x"0000",
    x"0D1D",
    x"1A16",
    x"26CA",
    x"3314",
    x"3ED5",
    x"49ED",
    x"543E",
    x"5DAC",
    x"661D",
    x"6D7C",
    x"73B3",
    x"78B3",
    x"7C6E",
    x"7ED9",
    x"7FEF",
    x"7FAC",
    x"7E11",
    x"7B23",
    x"76E9",
    x"716E",
    x"6AC2",
    x"62F7",
    x"5A21",
    x"5058",
    x"45B6",
    x"3A59",
    x"2E5F",
    x"21E7",
    x"1515",
    x"0809",
    x"FAE8",
    x"EDD5",
    x"E0F3",
    x"D464",
    x"C84B",
    x"BCC8",
    x"B1FA",
    x"A7FE",
    x"9EEF",
    x"96E5",
    x"8FF7",
    x"8A37",
    x"85B4",
    x"827A",
    x"8092",
    x"8002",
    x"80CB",
    x"82EA",
    x"865A",
    x"8B12",
    x"9105",
    x"9822",
    x"A058",
    x"A98F",
    x"B3AF",
    x"BE9D",
    x"CA3B",
    x"D66A",
    x"E308",
    x"EFF5",
    x"FD0D",
    x"0A2D",
    x"1732",
    x"23F8",
    x"305D",
    x"3C40",
    x"4780",
    x"5200",
    x"5BA3",
    x"644F",
    x"6BED",
    x"7269",
    x"77B0",
    x"7BB4",
    x"7E6C",
    x"7FCE",
    x"7FD9",
    x"7E8B",
    x"7BE8",
    x"77F8",
    x"72C4",
    x"6C5B",
    x"64CF",
    x"5C32",
    x"529E",
    x"482B",
    x"3CF5",
    x"311B",
    x"24BD",
    x"17FC",
    x"0AFA",
    x"FDDB",
    x"F0C2",
    x"E3D1",
    x"D72D",
    x"CAF6",
    x"BF4F",
    x"B455",
    x"AA28",
    x"A0E1",
    x"989B",
    x"916C",
    x"8B66",
    x"869B",
    x"8316",
    x"80E2",
    x"8005",
    x"8080",
    x"8252",
    x"8578",
    x"89E7",
    x"8F94",
    x"9670",
    x"9E69",
    x"A769",
    x"B157",
    x"BC19",
    x"C792",
    x"D3A3",
    x"E02B",
    x"ED09",
    x"FA1B",
    x"073C",
    x"144A",
    x"2121",
    x"2D9F",
    x"39A1",
    x"4509",
    x"4FB7",
    x"598E",
    x"6274",
    x"6A50",
    x"710E",
    x"769C",
    x"7AEA",
    x"7DED",
    x"7F9D",
    x"7FF5",
    x"7EF4",
    x"7C9D",
    x"78F7",
    x"740B",
    x"6DE6",
    x"6699",
    x"5E38",
    x"54D9",
    x"4A95",
    x"3F88",
    x"33D1",
    x"278E",
    x"1AE0",
    x"0DEA",
    x"00CE",
    x"F3B0",
    x"E6B3",
    x"D9FB",
    x"CDA9",
    x"C1DE",
    x"B6BB",
    x"AC5D",
    x"A2E1",
    x"9A5F",
    x"92EF",
    x"8CA5",
    x"8792",
    x"83C3",
    x"8143",
    x"8018",
    x"8046",
    x"81CC",
    x"84A6",
    x"88CC",
    x"8E33",
    x"94CD",
    x"9C87",
    x"A54E",
    x"AF09",
    x"B99D",
    x"C4F0",
    x"D0E2",
    x"DD52",
    x"EA20",
    x"F729",
    x"044A",
    x"115F",
    x"1E45",
    x"2ADA",
    x"36FC",
    x"4289",
    x"4D63",
    x"576C",
    x"608B",
    x"68A5",
    x"6FA5",
    x"7578",
    x"7A0F",
    x"7D5D",
    x"7F5A",
    x"7FFF",
    x"7F4B",
    x"7D41",
    x"79E5",
    x"7541",
    x"6F61",
    x"6855",
    x"6030",
    x"5708",
    x"4CF5",
    x"4213",
    x"3680",
    x"2A59",
    x"1DC0",
    x"10D7",
    x"03C1",
    x"F6A0",
    x"E999",
    x"DCCE",
    x"D062",
    x"C476",
    x"B92B",
    x"AE9E",
    x"A4ED",
    x"9C31",
    x"9482",
    x"8DF4",
    x"889A",
    x"8481",
    x"81B5",
    x"803D",
    x"801E",
    x"8157",
    x"83E5",
    x"87C1",
    x"8CE1",
    x"9338",
    x"9AB3",
    x"A33F",
    x"ACC5",
    x"B72C",
    x"C256",
    x"CE27",
    x"DA7E",
    x"E73A",
    x"F439",
    x"0157",
    x"0E72",
    x"1B66",
    x"2810",
    x"344E",
    x"3FFF",
    x"4B04",
    x"553F",
    x"5E94",
    x"66EB",
    x"6E2C",
    x"7444",
    x"7923",
    x"7CBC",
    x"7F05",
    x"7FF8",
    x"7F92",
    x"7DD4",
    x"7AC3",
    x"7668",
    x"70CE",
    x"6A03",
    x"621C",
    x"592C",
    x"4F4B",
    x"4495",
    x"3927",
    x"2D1E",
    x"209C",
    x"13C2",
    x"06B3",
    x"F992",
    x"EC82",
    x"DFA6",
    x"D322",
    x"C717",
    x"BBA5",
    x"B0EB",
    x"A706",
    x"9E10",
    x"9623",
    x"8F53",
    x"89B2",
    x"8550",
    x"8239",
    x"8074",
    x"8007",
    x"80F2",
    x"8334",
    x"86C6",
    x"8B9F",
    x"91B1",
    x"98EC",
    x"A13D",
    x"AA8E",
    x"B4C4",
    x"BFC5",
    x"CB73",
    x"D7AF",
    x"E457",
    x"F14A",
    x"FE64",
    x"0B83",
    x"1883",
    x"2540",
    x"319A",
    x"3D6D",
    x"489C",
    x"5306",
    x"5C91",
    x"6523",
    x"6CA4",
    x"7301",
    x"7827",
    x"7C0B",
    x"7E9F",
    x"7FDF",
    x"7FC7",
    x"7E56",
    x"7B91",
    x"777F",
    x"722B",
    x"6BA3",
    x"63FA",
    x"5B43",
    x"5196",
    x"470E",
    x"3BC6",
    x"2FDE",
    x"2374",
    x"16AB",
    x"09A4",
    x"FC84",
    x"EF6D",
    x"E283",
    x"D5E8",
    x"C9BF",
    x"BE27",
    x"B341",
    x"A92A",
    x"9FFD",
    x"97D3",
    x"90C1",
    x"8ADA",
    x"8630",
    x"82CD",
    x"80BC",
    x"8001",
    x"80A0",
    x"8295",
    x"85DC",
    x"8A6D",
    x"903A",
    x"9734",
    x"9F48",
    x"A861",
    x"B266",
    x"BD3D",
    x"C8C6",
    x"D4E5",
    x"E178",
    x"EE5D",
    x"FB72",
    x"0892",
    x"159C",
    x"226C",
    x"2EDF",
    x"3AD3",
    x"4629",
    x"50C2",
    x"5A82",
    x"634D",
    x"6B0E",
    x"71AE",
    x"771B",
    x"7B48",
    x"7E29",
    x"7FB5",
    x"7FEA",
    x"7EC6",
    x"7C4D",
    x"7885",
    x"7378",
    x"6D34",
    x"65CA",
    x"5D4E",
    x"53D7",
    x"497D",
    x"3E5E",
    x"3296",
    x"2647",
    x"1990",
    x"0C94",
    x"FF77",
    x"F25B",
    x"E563",
    x"D8B4",
    x"CC6E",
    x"C0B3",
    x"B5A3",
    x"AB5B",
    x"A1F7",
    x"9990",
    x"923D",
    x"8C12",
    x"8720",
    x"8372",
    x"8115",
    x"800D",
    x"805E",
    x"8207",
    x"8503",
    x"894A",
    x"8ED2",
    x"958A",
    x"9D61",
    x"A641",
    x"B013",
    x"BABD",
    x"C621",
    x"D221",
    x"DE9D",
    x"EB73",
    x"F880",
    x"05A1",
    x"12B3",
    x"1F92",
    x"2C1D",
    x"3831",
    x"43AD",
    x"4E73",
    x"5866",
    x"616A",
    x"6969",
    x"704B",
    x"75FF",
    x"7A75",
    x"7DA1",
    x"7F7A",
    x"7FFC",
    x"7F26",
    x"7CF9",
    x"797B",
    x"74B6",
    x"6EB7",
    x"678D",
    x"5F4C",
    x"560B",
    x"4BE2",
    x"40ED",
    x"3548",
    x"2914",
    x"1C72",
    x"0F83",
    x"026A",
    x"F54A",
    x"E848",
    x"DB85",
    x"CF24",
    x"C347",
    x"B80E",
    x"AD97",
    x"A3FD",
    x"9B5C",
    x"93C9",
    x"8D5A",
    x"8820",
    x"8429",
    x"817F",
    x"802A",
    x"802E",
    x"818A",
    x"843A",
    x"8838",
    x"8D79",
    x"93EE",
    x"9B86",
    x"A42D",
    x"ADCB",
    x"B847",
    x"C384",
    x"CF64",
    x"DBC7",
    x"E88B",
    x"F58F",
    x"02AE",
    x"0FC7",
    x"1CB5",
    x"2955",
    x"3587",
    x"4128",
    x"4C19",
    x"563E",
    x"5F7A",
    x"67B5",
    x"6ED9",
    x"74D2",
    x"7991",
    x"7D08",
    x"7F2E",
    x"7FFD",
    x"7F74",
    x"7D93",
    x"7A61",
    x"75E4",
    x"702A",
    x"6942",
    x"613E",
    x"5834",
    x"4E3D",
    x"4373",
    x"37F3",
    x"2BDC",
    x"1F50",
    x"126F",
    x"055C",
    x"F83B",
    x"EB2F",
    x"DE5B",
    x"D1E1",
    x"C5E4",
    x"BA83",
    x"AFDE",
    x"A610",
    x"9D35",
    x"9564",
    x"8EB2",
    x"8931",
    x"84F0",
    x"81FB",
    x"8059",
    x"800F",
    x"811E",
    x"8382",
    x"8736",
    x"8C30",
    x"9261",
    x"99B9",
    x"A225",
    x"AB8E",
    x"B5DB",
    x"C0EF",
    x"CCAD",
    x"D8F5",
    x"E5A6",
    x"F29F",
    x"FFBB",
    x"0CD9",
    x"19D3",
    x"2688",
    x"32D5",
    x"3E9A",
    x"49B5",
    x"540A",
    x"5D7D",
    x"65F4",
    x"6D58",
    x"7396",
    x"789C",
    x"7C5D",
    x"7ED0",
    x"7FED",
    x"7FB1",
    x"7E1D",
    x"7B35",
    x"7702",
    x"718E",
    x"6AE8",
    x"6322",
    x"5A51",
    x"508D",
    x"45F0",
    x"3A96",
    x"2E9F",
    x"222A",
    x"1559",
    x"084E",
    x"FB2D",
    x"EE19",
    x"E135",
    x"D4A5",
    x"C889",
    x"BD02",
    x"B230",
    x"A82F",
    x"9F1C",
    x"970D",
    x"9018",
    x"8A52",
    x"85C8",
    x"8287",
    x"8099",
    x"8002",
    x"80C3",
    x"82DB",
    x"8645",
    x"8AF6",
    x"90E3",
    x"97FA",
    x"A02B",
    x"A95D",
    x"B378",
    x"BE62",
    x"C9FD",
    x"D629",
    x"E2C6",
    x"EFB1",
    x"FCC9",
    x"09E9",
    x"16EE",
    x"23B6",
    x"301D",
    x"3C03",
    x"4747",
    x"51CB",
    x"5B73",
    x"6425",
    x"6BC8",
    x"724A",
    x"7797",
    x"7BA2",
    x"7E61",
    x"7FCB",
    x"7FDC",
    x"7E95",
    x"7BFA",
    x"7810",
    x"72E3",
    x"6C80",
    x"64F9",
    x"5C62",
    x"52D2",
    x"4863",
    x"3D31",
    x"315A",
    x"24FF",
    x"183F",
    x"0B3F",
    x"FE20",
    x"F106",
    x"E414",
    x"D76E",
    x"CB35",
    x"BF8A",
    x"B48D",
    x"AA5B",
    x"A10F",
    x"98C4",
    x"918E",
    x"8B83",
    x"86B0",
    x"8325",
    x"80EA",
    x"8006",
    x"807A",
    x"8245",
    x"8564",
    x"89CC",
    x"8F73",
    x"964A",
    x"9E3D",
    x"A737",
    x"B121",
    x"BBDF",
    x"C754",
    x"D362",
    x"DFE9",
    x"ECC6",
    x"F9D6",
    x"06F7",
    x"1406",
    x"20DE",
    x"2D5E",
    x"3964",
    x"44CF",
    x"4F81",
    x"595D",
    x"6248",
    x"6A2A",
    x"70EE",
    x"7682",
    x"7AD7",
    x"7DE1",
    x"7F97",
    x"7FF6",
    x"7EFD",
    x"7CAD",
    x"790D",
    x"7428",
    x"6E09",
    x"66C2",
    x"5E66",
    x"550C",
    x"4ACD",
    x"3FC4",
    x"3410",
    x"27CF",
    x"1B23",
    x"0E2E",
    x"0113",
    x"F3F4",
    x"E6F7",
    x"DA3C",
    x"CDE8",
    x"C21A",
    x"B6F3",
    x"AC91",
    x"A310",
    x"9A89",
    x"9313",
    x"8CC3",
    x"87A9",
    x"83D4",
    x"814D",
    x"801B",
    x"8042",
    x"81C0",
    x"8493",
    x"88B3",
    x"8E14",
    x"94A7",
    x"9C5C",
    x"A51D",
    x"AED3",
    x"B964",
    x"C4B3",
    x"D0A2",
    x"DD10",
    x"E9DD",
    x"F6E5",
    x"0405",
    x"111B",
    x"1E03",
    x"2A99",
    x"36BE",
    x"424E",
    x"4D2C",
    x"573A",
    x"605D",
    x"687D",
    x"6F83",
    x"755D",
    x"79FA",
    x"7D4F",
    x"7F53",
    x"7FFF",
    x"7F53",
    x"7D4F",
    x"79FA",
    x"755D",
    x"6F83",
    x"687D",
    x"605D",
    x"573A",
    x"4D2C",
    x"424E",
    x"36BE",
    x"2A99",
    x"1E03",
    x"111B",
    x"0405",
    x"F6E5",
    x"E9DD",
    x"DD10",
    x"D0A2",
    x"C4B3",
    x"B964",
    x"AED3",
    x"A51D",
    x"9C5C",
    x"94A7",
    x"8E14",
    x"88B3",
    x"8493",
    x"81C0",
    x"8042",
    x"801B",
    x"814D",
    x"83D4",
    x"87A9",
    x"8CC3",
    x"9313",
    x"9A89",
    x"A310",
    x"AC91",
    x"B6F3",
    x"C21A",
    x"CDE8",
    x"DA3C",
    x"E6F7",
    x"F3F4",
    x"0113",
    x"0E2E",
    x"1B23",
    x"27CF",
    x"3410",
    x"3FC4",
    x"4ACD",
    x"550C",
    x"5E66",
    x"66C2",
    x"6E09",
    x"7428",
    x"790D",
    x"7CAD",
    x"7EFD",
    x"7FF6",
    x"7F97",
    x"7DE1",
    x"7AD7",
    x"7682",
    x"70EE",
    x"6A2A",
    x"6248",
    x"595D",
    x"4F81",
    x"44CF",
    x"3964",
    x"2D5E",
    x"20DE",
    x"1406",
    x"06F7",
    x"F9D6",
    x"ECC6",
    x"DFE9",
    x"D362",
    x"C754",
    x"BBDF",
    x"B121",
    x"A737",
    x"9E3D",
    x"964A",
    x"8F73",
    x"89CC",
    x"8564",
    x"8245",
    x"807A",
    x"8006",
    x"80EA",
    x"8325",
    x"86B0",
    x"8B83",
    x"918E",
    x"98C4",
    x"A10F",
    x"AA5B",
    x"B48D",
    x"BF8A",
    x"CB35",
    x"D76E",
    x"E414",
    x"F106",
    x"FE20",
    x"0B3F",
    x"183F",
    x"24FF",
    x"315A",
    x"3D31",
    x"4863",
    x"52D2",
    x"5C62",
    x"64F9",
    x"6C80",
    x"72E3",
    x"7810",
    x"7BFA",
    x"7E95",
    x"7FDC",
    x"7FCB",
    x"7E61",
    x"7BA2",
    x"7797",
    x"724A",
    x"6BC8",
    x"6425",
    x"5B73",
    x"51CB",
    x"4747",
    x"3C03",
    x"301D",
    x"23B6",
    x"16EE",
    x"09E9",
    x"FCC9",
    x"EFB1",
    x"E2C6",
    x"D629",
    x"C9FD",
    x"BE62",
    x"B378",
    x"A95D",
    x"A02B",
    x"97FA",
    x"90E3",
    x"8AF6",
    x"8645",
    x"82DB",
    x"80C3",
    x"8002",
    x"8099",
    x"8287",
    x"85C8",
    x"8A52",
    x"9018",
    x"970D",
    x"9F1C",
    x"A82F",
    x"B230",
    x"BD02",
    x"C889",
    x"D4A5",
    x"E135",
    x"EE19",
    x"FB2D",
    x"084E",
    x"1559",
    x"222A",
    x"2E9F",
    x"3A96",
    x"45F0",
    x"508D",
    x"5A51",
    x"6322",
    x"6AE8",
    x"718E",
    x"7702",
    x"7B35",
    x"7E1D",
    x"7FB1",
    x"7FED",
    x"7ED0",
    x"7C5D",
    x"789C",
    x"7396",
    x"6D58",
    x"65F4",
    x"5D7D",
    x"540A",
    x"49B5",
    x"3E9A",
    x"32D5",
    x"2688",
    x"19D3",
    x"0CD9",
    x"FFBB",
    x"F29F",
    x"E5A6",
    x"D8F5",
    x"CCAD",
    x"C0EF",
    x"B5DB",
    x"AB8E",
    x"A225",
    x"99B9",
    x"9261",
    x"8C30",
    x"8736",
    x"8382",
    x"811E",
    x"800F",
    x"8059",
    x"81FB",
    x"84F0",
    x"8931",
    x"8EB2",
    x"9564",
    x"9D35",
    x"A610",
    x"AFDE",
    x"BA83",
    x"C5E4",
    x"D1E1",
    x"DE5B",
    x"EB2F",
    x"F83B",
    x"055C",
    x"126F",
    x"1F50",
    x"2BDC",
    x"37F3",
    x"4373",
    x"4E3D",
    x"5834",
    x"613E",
    x"6942",
    x"702A",
    x"75E4",
    x"7A61",
    x"7D93",
    x"7F74",
    x"7FFD",
    x"7F2E",
    x"7D08",
    x"7991",
    x"74D2",
    x"6ED9",
    x"67B5",
    x"5F7A",
    x"563E",
    x"4C19",
    x"4128",
    x"3587",
    x"2955",
    x"1CB5",
    x"0FC7",
    x"02AE",
    x"F58F",
    x"E88B",
    x"DBC7",
    x"CF64",
    x"C384",
    x"B847",
    x"ADCB",
    x"A42D",
    x"9B86",
    x"93EE",
    x"8D79",
    x"8838",
    x"843A",
    -- nota 08
    x"0000",
    x"0DE4",
    x"1B9D",
    x"2903",
    x"35ED",
    x"4235",
    x"4DB3",
    x"5847",
    x"61D1",
    x"6A32",
    x"7152",
    x"771C",
    x"7B7E",
    x"7E6A",
    x"7FD8",
    x"7FC4",
    x"7E2D",
    x"7B19",
    x"7691",
    x"70A2",
    x"695F",
    x"60DD",
    x"5737",
    x"4C88",
    x"40F3",
    x"3499",
    x"27A0",
    x"1A2F",
    x"0C6F",
    x"FE89",
    x"F0A8",
    x"E2F5",
    x"D59A",
    x"C8C0",
    x"BC8C",
    x"B124",
    x"A6AB",
    x"9D3F",
    x"94FF",
    x"8E01",
    x"885D",
    x"8422",
    x"815D",
    x"8018",
    x"8055",
    x"8214",
    x"8550",
    x"89FE",
    x"9012",
    x"9778",
    x"A019",
    x"A9DD",
    x"B4A6",
    x"C052",
    x"CCBE",
    x"D9C6",
    x"E741",
    x"F507",
    x"02EE",
    x"10CC",
    x"1E77",
    x"2BC7",
    x"3892",
    x"44B2",
    x"5002",
    x"5A60",
    x"63AE",
    x"6BCD",
    x"72A7",
    x"7827",
    x"7C3B",
    x"7ED7",
    x"7FF4",
    x"7F8E",
    x"7DA7",
    x"7A43",
    x"756F",
    x"6F37",
    x"67AE",
    x"5EED",
    x"550C",
    x"4A2A",
    x"3E68",
    x"31EA",
    x"24D4",
    x"174F",
    x"0984",
    x"FB9C",
    x"EDC1",
    x"E01D",
    x"D2DA",
    x"C61F",
    x"BA13",
    x"AEDB",
    x"A498",
    x"9B69",
    x"936A",
    x"8CB4",
    x"875A",
    x"836D",
    x"80F9",
    x"8004",
    x"8093",
    x"82A3",
    x"862D",
    x"8B29",
    x"9185",
    x"992F",
    x"A210",
    x"AC0E",
    x"B709",
    x"C2E0",
    x"CF70",
    x"DC94",
    x"EA22",
    x"F7F2",
    x"05DB",
    x"13B2",
    x"214D",
    x"2E84",
    x"3B2E",
    x"4726",
    x"5246",
    x"5C6D",
    x"657D",
    x"6D5A",
    x"73ED",
    x"7921",
    x"7CE7",
    x"7F33",
    x"7FFF",
    x"7F48",
    x"7D10",
    x"795D",
    x"743C",
    x"6DBC",
    x"65F0",
    x"5CEF",
    x"52D6",
    x"47C2",
    x"3BD5",
    x"2F34",
    x"2204",
    x"146C",
    x"0697",
    x"F8AF",
    x"EADC",
    x"DD49",
    x"D01F",
    x"C386",
    x"B7A4",
    x"AC9C",
    x"A291",
    x"99A0",
    x"91E5",
    x"8B76",
    x"8668",
    x"82C9",
    x"80A5",
    x"8002",
    x"80E2",
    x"8342",
    x"871C",
    x"8C62",
    x"9307",
    x"9AF5",
    x"A414",
    x"AE49",
    x"B975",
    x"C577",
    x"D229",
    x"DF66",
    x"ED06",
    x"FADF",
    x"08C7",
    x"1695",
    x"241F",
    x"313C",
    x"3DC3",
    x"4990",
    x"547F",
    x"5E6E",
    x"673F",
    x"6ED9",
    x"7523",
    x"7A0B",
    x"7D82",
    x"7F7E",
    x"7FF8",
    x"7EF0",
    x"7C68",
    x"7867",
    x"72FB",
    x"6C33",
    x"6424",
    x"5AE6",
    x"5095",
    x"4551",
    x"393B",
    x"2C78",
    x"1F2F",
    x"1187",
    x"03AA",
    x"F5C3",
    x"E7FA",
    x"DA7A",
    x"CD6B",
    x"C0F6",
    x"B53E",
    x"AA69",
    x"A097",
    x"97E5",
    x"906E",
    x"8A48",
    x"8586",
    x"8236",
    x"8063",
    x"8011",
    x"8142",
    x"83F3",
    x"881A",
    x"8DAC",
    x"9497",
    x"9CC8",
    x"A624",
    x"B090",
    x"BBEC",
    x"C816",
    x"D4E8",
    x"E23E",
    x"EFED",
    x"FDCC",
    x"0BB3",
    x"1976",
    x"26EC",
    x"33EC",
    x"4050",
    x"4BF1",
    x"56AC",
    x"6061",
    x"68F3",
    x"7048",
    x"7649",
    x"7AE5",
    x"7E0D",
    x"7FB8",
    x"7FE1",
    x"7E87",
    x"7BAF",
    x"7761",
    x"71AA",
    x"6A9B",
    x"624A",
    x"58D0",
    x"4E49",
    x"42D6",
    x"3698",
    x"29B6",
    x"1C55",
    x"0E9F",
    x"00BD",
    x"F2D8",
    x"E51B",
    x"D7B0",
    x"CABE",
    x"BE6D",
    x"B2E3",
    x"A842",
    x"9EAA",
    x"9638",
    x"8F06",
    x"8929",
    x"84B4",
    x"81B4",
    x"8031",
    x"8031",
    x"81B4",
    x"84B4",
    x"8929",
    x"8F05",
    x"9636",
    x"9EA8",
    x"A840",
    x"B2E1",
    x"BE6B",
    x"CABC",
    x"D7AD",
    x"E519",
    x"F2D6",
    x"00BA",
    x"0E9D",
    x"1C53",
    x"29B3",
    x"3696",
    x"42D4",
    x"4E47",
    x"58CE",
    x"6248",
    x"6A99",
    x"71A8",
    x"7760",
    x"7BAE",
    x"7E87",
    x"7FE1",
    x"7FB8",
    x"7E0D",
    x"7AE6",
    x"764A",
    x"7049",
    x"68F5",
    x"6063",
    x"56AE",
    x"4BF3",
    x"4052",
    x"33EF",
    x"26EE",
    x"1978",
    x"0BB5",
    x"FDCF",
    x"EFEF",
    x"E240",
    x"D4EB",
    x"C818",
    x"BBEE",
    x"B092",
    x"A626",
    x"9CC9",
    x"9499",
    x"8DAD",
    x"881B",
    x"83F3",
    x"8143",
    x"8011",
    x"8063",
    x"8236",
    x"8585",
    x"8A47",
    x"906D",
    x"97E3",
    x"A095",
    x"AA67",
    x"B53C",
    x"C0F3",
    x"CD69",
    x"DA77",
    x"E7F7",
    x"F5C0",
    x"03A8",
    x"1184",
    x"1F2C",
    x"2C75",
    x"3938",
    x"454E",
    x"5093",
    x"5AE4",
    x"6422",
    x"6C31",
    x"72FA",
    x"7866",
    x"7C67",
    x"7EF0",
    x"7FF8",
    x"7F7E",
    x"7D83",
    x"7A0C",
    x"7524",
    x"6EDA",
    x"6741",
    x"5E6F",
    x"5481",
    x"4992",
    x"3DC5",
    x"313E",
    x"2422",
    x"1698",
    x"08CA",
    x"FAE2",
    x"ED09",
    x"DF69",
    x"D22C",
    x"C579",
    x"B978",
    x"AE4B",
    x"A416",
    x"9AF6",
    x"9308",
    x"8C64",
    x"871D",
    x"8343",
    x"80E2",
    x"8002",
    x"80A5",
    x"82C9",
    x"8667",
    x"8B75",
    x"91E3",
    x"999F",
    x"A28F",
    x"AC9A",
    x"B7A2",
    x"C384",
    x"D01D",
    x"DD47",
    x"EAD9",
    x"F8AC",
    x"0695",
    x"146A",
    x"2201",
    x"2F31",
    x"3BD3",
    x"47C0",
    x"52D4",
    x"5CEE",
    x"65EE",
    x"6DBB",
    x"743B",
    x"795D",
    x"7D0F",
    x"7F47",
    x"7FFF",
    x"7F33",
    x"7CE7",
    x"7922",
    x"73EE",
    x"6D5C",
    x"657F",
    x"5C6F",
    x"5248",
    x"4728",
    x"3B31",
    x"2E87",
    x"2150",
    x"13B5",
    x"05DE",
    x"F7F5",
    x"EA24",
    x"DC96",
    x"CF73",
    x"C2E2",
    x"B70B",
    x"AC10",
    x"A212",
    x"9931",
    x"9186",
    x"8B2A",
    x"862E",
    x"82A3",
    x"8093",
    x"8004",
    x"80F8",
    x"836D",
    x"8759",
    x"8CB3",
    x"9369",
    x"9B67",
    x"A496",
    x"AED9",
    x"BA11",
    x"C61D",
    x"D2D7",
    x"E01B",
    x"EDBE",
    x"FB99",
    x"0981",
    x"174D",
    x"24D2",
    x"31E7",
    x"3E66",
    x"4A28",
    x"550A",
    x"5EEB",
    x"67AD",
    x"6F35",
    x"756D",
    x"7A43",
    x"7DA6",
    x"7F8E",
    x"7FF4",
    x"7ED7",
    x"7C3B",
    x"7827",
    x"72A8",
    x"6BCF",
    x"63AF",
    x"5A62",
    x"5004",
    x"44B4",
    x"3894",
    x"2BC9",
    x"1E7A",
    x"10CE",
    x"02F0",
    x"F509",
    x"E743",
    x"D9C8",
    x"CCC0",
    x"C054",
    x"B4A8",
    x"A9DF",
    x"A01B",
    x"9779",
    x"9013",
    x"89FF",
    x"8550",
    x"8214",
    x"8055",
    x"8018",
    x"815D",
    x"8421",
    x"885C",
    x"8E00",
    x"94FD",
    x"9D3E",
    x"A6A9",
    x"B122",
    x"BC8A",
    x"C8BD",
    x"D598",
    x"E2F3",
    x"F0A5",
    x"FE87",
    x"0C6C",
    x"1A2C",
    x"279D",
    x"3496",
    x"40F0",
    x"4C86",
    x"5735",
    x"60DB",
    x"695D",
    x"70A1",
    x"7690",
    x"7B18",
    x"7E2D",
    x"7FC4",
    x"7FD8",
    x"7E6B",
    x"7B7E",
    x"771D",
    x"7154",
    x"6A33",
    x"61D2",
    x"5849",
    x"4DB5",
    x"4237",
    x"35F0",
    x"2906",
    x"1BA0",
    x"0DE6",
    x"0003",
    x"F21F",
    x"E465",
    x"D6FF",
    x"CA15",
    x"BDCE",
    x"B24F",
    x"A7BA",
    x"9E31",
    x"95CF",
    x"8EAF",
    x"88E5",
    x"8483",
    x"8196",
    x"8028",
    x"803C",
    x"81D2",
    x"84E6",
    x"896E",
    x"8F5D",
    x"96A0",
    x"9F21",
    x"A8C8",
    x"B376",
    x"BF0B",
    x"CB65",
    x"D85E",
    x"E5CF",
    x"F38F",
    x"0174",
    x"0F55",
    x"1D08",
    x"2A63",
    x"373E",
    x"4372",
    x"4EDA",
    x"5954",
    x"62BF",
    x"6B00",
    x"71FE",
    x"77A2",
    x"7BDE",
    x"7EA2",
    x"7FE8",
    x"7FAB",
    x"7DED",
    x"7AB1",
    x"7603",
    x"6FEF",
    x"688A",
    x"5FE8",
    x"5625",
    x"4B5D",
    x"3FB1",
    x"3344",
    x"263D",
    x"18C2",
    x"0AFC",
    x"FD15",
    x"EF37",
    x"E18B",
    x"D43C",
    x"C771",
    x"BB50",
    x"B000",
    x"A5A1",
    x"9C54",
    x"9434",
    x"8D5A",
    x"87DA",
    x"83C6",
    x"8129",
    x"800C",
    x"8071",
    x"8259",
    x"85BC",
    x"8A90",
    x"90C8",
    x"9850",
    x"A112",
    x"AAF2",
    x"B5D4",
    x"C196",
    x"CE14",
    x"DB2A",
    x"E8AE",
    x"F67A",
    x"0462",
    x"123D",
    x"1FE0",
    x"2D24",
    x"39DF",
    x"45EB",
    x"5123",
    x"5B67",
    x"6495",
    x"6C94",
    x"734B",
    x"78A5",
    x"7C92",
    x"7F07",
    x"7FFC",
    x"7F6D",
    x"7D5E",
    x"79D3",
    x"74D8",
    x"6E7C",
    x"66D2",
    x"5DF1",
    x"53F4",
    x"48FA",
    x"3D22",
    x"3092",
    x"236F",
    x"15E1",
    x"0810",
    x"FA28",
    x"EC51",
    x"DEB5",
    x"D17E",
    x"C4D4",
    x"B8DC",
    x"ADBC",
    x"A395",
    x"9A84",
    x"92A7",
    x"8C14",
    x"86E0",
    x"831A",
    x"80CD",
    x"8001",
    x"80B8",
    x"82F0",
    x"86A2",
    x"8BC3",
    x"9243",
    x"9A0F",
    x"A30F",
    x"AD28",
    x"B83C",
    x"C428",
    x"D0CA",
    x"DDFA",
    x"EB91",
    x"F966",
    x"074F",
    x"1522",
    x"22B4",
    x"2FDE",
    x"3C78",
    x"485A",
    x"5362",
    x"5D6D",
    x"665E",
    x"6E1A",
    x"7489",
    x"7997",
    x"7D36",
    x"7F5B",
    x"7FFE",
    x"7F1E",
    x"7CBE",
    x"78E5",
    x"739F",
    x"6CFA",
    x"650D",
    x"5BEE",
    x"51B9",
    x"468D",
    x"3A8B",
    x"2DD9",
    x"209C",
    x"12FD",
    x"0524",
    x"F73B",
    x"E96D",
    x"DBE3",
    x"CEC7",
    x"C23F",
    x"B672",
    x"AB83",
    x"A194",
    x"98C2",
    x"9129",
    x"8ADE",
    x"85F6",
    x"827E",
    x"8082",
    x"8008",
    x"8110",
    x"8398",
    x"8798",
    x"8D04",
    x"93CC",
    x"9BDB",
    x"A519",
    x"AF69",
    x"BAAD",
    x"C6C3",
    x"D386",
    x"E0CF",
    x"EE77",
    x"FC53",
    x"0A3B",
    x"1804",
    x"2584",
    x"3292",
    x"3F08",
    x"4AC0",
    x"5595",
    x"5F67",
    x"681A",
    x"6F91",
    x"75B7",
    x"7A79",
    x"7DC9",
    x"7F9D",
    x"7FEF",
    x"7EBE",
    x"7C0E",
    x"77E7",
    x"7255",
    x"6B6A",
    x"633A",
    x"59DE",
    x"4F72",
    x"4417",
    x"37ED",
    x"2B1A",
    x"1DC5",
    x"1016",
    x"0236",
    x"F450",
    x"E68D",
    x"D917",
    x"CC16",
    x"BFB3",
    x"B411",
    x"A956",
    x"9FA0",
    x"970E",
    x"8FB9",
    x"89B8",
    x"851C",
    x"81F3",
    x"8048",
    x"801F",
    x"8178",
    x"8450",
    x"889E",
    x"8E55",
    x"9564",
    x"9DB4",
    x"A72E",
    x"B1B5",
    x"BD28",
    x"C965",
    x"D648",
    x"E3A8",
    x"F15E",
    x"FF41",
    x"0D25",
    x"1AE2",
    x"284E",
    x"3540",
    x"4190",
    x"4D1B",
    x"57BD",
    x"6155",
    x"69C7",
    x"70F9",
    x"76D6",
    x"7B4B",
    x"7E4C",
    x"7FCE",
    x"7FCF",
    x"7E4D",
    x"7B4D",
    x"76D8",
    x"70FD",
    x"69CB",
    x"615A",
    x"57C2",
    x"4D21",
    x"4197",
    x"3547",
    x"2855",
    x"1AEA",
    x"0D2D",
    x"FF48",
    x"F166",
    x"E3B0",
    x"D64F",
    x"C96C",
    x"BD2F",
    x"B1BB",
    x"A734",
    x"9DB9",
    x"9568",
    x"8E59",
    x"88A1",
    x"8452",
    x"817A",
    x"801F",
    x"8048",
    x"81F2",
    x"851A",
    x"89B5",
    x"8FB5",
    x"970A",
    x"9F9B",
    x"A950",
    x"B40B",
    x"BFAC",
    x"CC0F",
    x"D90F",
    x"E685",
    x"F448",
    x"022E",
    x"100E",
    x"1DBD",
    x"2B13",
    x"37E6",
    x"4410",
    x"4F6C",
    x"59D9",
    x"6335",
    x"6B66",
    x"7252",
    x"77E4",
    x"7C0C",
    x"7EBD",
    x"7FEF",
    x"7F9E",
    x"7DCB",
    x"7A7C",
    x"75BA",
    x"6F95",
    x"681E",
    x"5F6D",
    x"559B",
    x"4AC6",
    x"3F0F",
    x"3299",
    x"258B",
    x"180B",
    x"0A42",
    x"FC5B",
    x"EE7E",
    x"E0D6",
    x"D38D",
    x"C6CA",
    x"BAB4",
    x"AF6F",
    x"A51E",
    x"9BE0",
    x"93D0",
    x"8D08",
    x"879B",
    x"839A",
    x"8111",
    x"8008",
    x"8081",
    x"827D",
    x"85F3",
    x"8ADB",
    x"9125",
    x"98BE",
    x"A18F",
    x"AB7E",
    x"B66C",
    x"C238",
    x"CEC0",
    x"DBDC",
    x"E966",
    x"F733",
    x"051C",
    x"12F5",
    x"2095",
    x"2DD2",
    x"3A85",
    x"4686",
    x"51B3",
    x"5BE8",
    x"6508",
    x"6CF6",
    x"739B",
    x"78E3",
    x"7CBD",
    x"7F1D",
    x"7FFE",
    x"7F5B",
    x"7D38",
    x"799A",
    x"748C",
    x"6E1E",
    x"6663",
    x"5D72",
    x"5367",
    x"4860",
    x"3C7E",
    x"2FE5",
    x"22BC",
    x"1529",
    x"0756",
    x"F96E",
    x"EB99",
    x"DE01",
    x"D0D1",
    x"C42F",
    x"B842",
    x"AD2E",
    x"A314",
    x"9A13",
    x"9247",
    x"8BC6",
    x"86A4",
    x"82F2",
    x"80B9",
    x"8001",
    x"80CC",
    x"8318",
    x"86DD",
    x"8C11",
    x"92A3",
    x"9A80",
    x"A38F",
    x"ADB6",
    x"B8D6",
    x"C4CD",
    x"D177",
    x"DEAE",
    x"EC49",
    x"FA20",
    x"0809",
    x"15D9",
    x"2367",
    x"308B",
    x"3D1B",
    x"48F3",
    x"53EF",
    x"5DEC",
    x"66CE",
    x"6E78",
    x"74D5",
    x"79D1",
    x"7D5C",
    x"7F6D",
    x"7FFC",
    x"7F08",
    x"7C94",
    x"78A8",
    x"734E",
    x"6C98",
    x"649A",
    x"5B6C",
    x"5129",
    x"45F1",
    x"39E6",
    x"2D2B",
    x"1FE8",
    x"1244",
    x"046A",
    x"F681",
    x"E8B6",
    x"DB31",
    x"CE1B",
    x"C19C",
    x"B5DA",
    x"AAF8",
    x"A117",
    x"9855",
    x"90CC",
    x"8A94",
    x"85BE",
    -- nota 09
    x"0000",
    x"0EB6",
    x"1D3A",
    x"2B5B",
    x"38E9",
    x"45B6",
    x"5196",
    x"5C62",
    x"65F4",
    x"6E2C",
    x"74EE",
    x"7A24",
    x"7DBB",
    x"7FA7",
    x"7FE2",
    x"7E6C",
    x"7B48",
    x"7682",
    x"702A",
    x"6855",
    x"5F1F",
    x"54A5",
    x"490D",
    x"3C7C",
    x"2F1E",
    x"2121",
    x"12B3",
    x"0405",
    x"F54A",
    x"E6B3",
    x"D872",
    x"CAB8",
    x"BDB2",
    x"B18D",
    x"A672",
    x"9C87",
    x"93EE",
    x"8CC3",
    x"8720",
    x"8316",
    x"80B5",
    x"8003",
    x"8103",
    x"83B3",
    x"8808",
    x"8DF4",
    x"9564",
    x"9E3D",
    x"A861",
    x"B3AF",
    x"C001",
    x"CD2B",
    x"DB01",
    x"E955",
    x"F7F7",
    x"06B3",
    x"1559",
    x"23B6",
    x"319A",
    x"3ED5",
    x"4B3C",
    x"56A3",
    x"60E4",
    x"69DD",
    x"716E",
    x"777F",
    x"7BFA",
    x"7ED0",
    x"7FF8",
    x"7F6E",
    x"7D33",
    x"7950",
    x"73D0",
    x"6CC8",
    x"644F",
    x"5A82",
    x"4F81",
    x"4373",
    x"3680",
    x"28D3",
    x"1A9D",
    x"0C0C",
    x"FD52",
    x"EEA1",
    x"E02B",
    x"D221",
    x"C4B3",
    x"B80E",
    x"AC5D",
    x"A1C8",
    x"9873",
    x"907D",
    x"8A01",
    x"8516",
    x"81CC",
    x"802E",
    x"8042",
    x"8207",
    x"8578",
    x"8A88",
    x"9127",
    x"993E",
    x"A2B2",
    x"AD62",
    x"B92B",
    x"C5E4",
    x"D362",
    x"E178",
    x"EFF5",
    x"FEA9",
    x"0D61",
    x"1BEC",
    x"2A18",
    x"37B5",
    x"4495",
    x"508D",
    x"5B73",
    x"6523",
    x"6D7C",
    x"7461",
    x"79BB",
    x"7D79",
    x"7F8C",
    x"7FEF",
    x"7E9F",
    x"7BA2",
    x"7702",
    x"70CE",
    x"691B",
    x"6003",
    x"55A5",
    x"4A25",
    x"3DAA",
    x"305D",
    x"226C",
    x"1406",
    x"055C",
    x"F6A0",
    x"E804",
    x"D9B9",
    x"CBF0",
    x"BED8",
    x"B29D",
    x"A769",
    x"9D61",
    x"94A7",
    x"8D5A",
    x"8792",
    x"8363",
    x"80DA",
    x"8001",
    x"80DA",
    x"8363",
    x"8792",
    x"8D5A",
    x"94A7",
    x"9D61",
    x"A769",
    x"B29D",
    x"BED8",
    x"CBF0",
    x"D9B9",
    x"E804",
    x"F6A0",
    x"055C",
    x"1406",
    x"226C",
    x"305D",
    x"3DAA",
    x"4A25",
    x"55A5",
    x"6003",
    x"691B",
    x"70CE",
    x"7702",
    x"7BA2",
    x"7E9F",
    x"7FEF",
    x"7F8C",
    x"7D79",
    x"79BB",
    x"7461",
    x"6D7C",
    x"6523",
    x"5B73",
    x"508D",
    x"4495",
    x"37B5",
    x"2A18",
    x"1BEC",
    x"0D61",
    x"FEA9",
    x"EFF5",
    x"E178",
    x"D362",
    x"C5E4",
    x"B92B",
    x"AD62",
    x"A2B2",
    x"993E",
    x"9127",
    x"8A88",
    x"8578",
    x"8207",
    x"8042",
    x"802E",
    x"81CC",
    x"8516",
    x"8A01",
    x"907D",
    x"9873",
    x"A1C8",
    x"AC5D",
    x"B80E",
    x"C4B3",
    x"D221",
    x"E02B",
    x"EEA1",
    x"FD52",
    x"0C0C",
    x"1A9D",
    x"28D3",
    x"3680",
    x"4373",
    x"4F81",
    x"5A82",
    x"644F",
    x"6CC8",
    x"73D0",
    x"7950",
    x"7D33",
    x"7F6E",
    x"7FF8",
    x"7ED0",
    x"7BFA",
    x"777F",
    x"716E",
    x"69DD",
    x"60E4",
    x"56A3",
    x"4B3C",
    x"3ED5",
    x"319A",
    x"23B6",
    x"1559",
    x"06B3",
    x"F7F7",
    x"E955",
    x"DB01",
    x"CD2B",
    x"C000",
    x"B3AF",
    x"A861",
    x"9E3D",
    x"9564",
    x"8DF4",
    x"8808",
    x"83B3",
    x"8103",
    x"8003",
    x"80B5",
    x"8316",
    x"8720",
    x"8CC3",
    x"93EE",
    x"9C87",
    x"A672",
    x"B18D",
    x"BDB2",
    x"CAB8",
    x"D872",
    x"E6B3",
    x"F54A",
    x"0405",
    x"12B3",
    x"2121",
    x"2F1E",
    x"3C7C",
    x"490D",
    x"54A5",
    x"5F1F",
    x"6855",
    x"702A",
    x"7682",
    x"7B48",
    x"7E6C",
    x"7FE2",
    x"7FA7",
    x"7DBB",
    x"7A24",
    x"74EE",
    x"6E2C",
    x"65F4",
    x"5C62",
    x"5196",
    x"45B6",
    x"38E9",
    x"2B5B",
    x"1D3A",
    x"0EB6",
    x"0000",
    x"F14A",
    x"E2C6",
    x"D4A5",
    x"C717",
    x"BA4A",
    x"AE6A",
    x"A39E",
    x"9A0C",
    x"91D4",
    x"8B12",
    x"85DC",
    x"8245",
    x"8059",
    x"801E",
    x"8194",
    x"84B8",
    x"897E",
    x"8FD6",
    x"97AB",
    x"A0E1",
    x"AB5B",
    x"B6F3",
    x"C384",
    x"D0E2",
    x"DEDF",
    x"ED4D",
    x"FBFB",
    x"0AB6",
    x"194D",
    x"278E",
    x"3548",
    x"424E",
    x"4E73",
    x"598E",
    x"6379",
    x"6C12",
    x"733D",
    x"78E0",
    x"7CEA",
    x"7F4B",
    x"7FFD",
    x"7EFD",
    x"7C4D",
    x"77F8",
    x"720C",
    x"6A9C",
    x"61C3",
    x"579F",
    x"4C51",
    x"4000",
    x"32D5",
    x"24FF",
    x"16AB",
    x"0809",
    x"F94D",
    x"EAA7",
    x"DC4A",
    x"CE66",
    x"C12B",
    x"B4C4",
    x"A95D",
    x"9F1C",
    x"9623",
    x"8E92",
    x"8881",
    x"8406",
    x"8130",
    x"8008",
    x"8092",
    x"82CD",
    x"86B0",
    x"8C30",
    x"9338",
    x"9BB1",
    x"A57E",
    x"B07F",
    x"BC8D",
    x"C980",
    x"D72D",
    x"E563",
    x"F3F4",
    x"02AE",
    x"115F",
    x"1FD5",
    x"2DDF",
    x"3B4D",
    x"47F2",
    x"53A3",
    x"5E38",
    x"678D",
    x"6F83",
    x"75FF",
    x"7AEA",
    x"7E34",
    x"7FD2",
    x"7FBE",
    x"7DF9",
    x"7A88",
    x"7578",
    x"6ED9",
    x"66C2",
    x"5D4E",
    x"529E",
    x"46D5",
    x"3A1C",
    x"2C9E",
    x"1E88",
    x"100B",
    x"0157",
    x"F29F",
    x"E414",
    x"D5E8",
    x"C84B",
    x"BB6B",
    x"AF73",
    x"A48D",
    x"9ADD",
    x"9284",
    x"8B9F",
    x"8645",
    x"8287",
    x"8074",
    x"8011",
    x"8161",
    x"845E",
    x"88FE",
    x"8F32",
    x"96E5",
    x"9FFD",
    x"AA5B",
    x"B5DB",
    x"C256",
    x"CFA3",
    x"DD94",
    x"EBFA",
    x"FAA4",
    x"0960",
    x"17FC",
    x"2647",
    x"3410",
    x"4128",
    x"4D63",
    x"5897",
    x"629F",
    x"6B59",
    x"72A6",
    x"786E",
    x"7C9D",
    x"7F26",
    x"7FFF",
    x"7F26",
    x"7C9D",
    x"786E",
    x"72A6",
    x"6B59",
    x"629F",
    x"5897",
    x"4D63",
    x"4128",
    x"3410",
    x"2647",
    x"17FC",
    x"0960",
    x"FAA4",
    x"EBFA",
    x"DD94",
    x"CFA3",
    x"C256",
    x"B5DB",
    x"AA5B",
    x"9FFD",
    x"96E5",
    x"8F32",
    x"88FE",
    x"845E",
    x"8161",
    x"8011",
    x"8074",
    x"8287",
    x"8645",
    x"8B9F",
    x"9284",
    x"9ADD",
    x"A48D",
    x"AF73",
    x"BB6B",
    x"C84B",
    x"D5E8",
    x"E414",
    x"F29F",
    x"0157",
    x"100B",
    x"1E88",
    x"2C9E",
    x"3A1C",
    x"46D5",
    x"529E",
    x"5D4E",
    x"66C2",
    x"6ED9",
    x"7578",
    x"7A88",
    x"7DF9",
    x"7FBE",
    x"7FD2",
    x"7E34",
    x"7AEA",
    x"75FF",
    x"6F83",
    x"678D",
    x"5E38",
    x"53A3",
    x"47F2",
    x"3B4D",
    x"2DDF",
    x"1FD5",
    x"115F",
    x"02AE",
    x"F3F4",
    x"E563",
    x"D72D",
    x"C980",
    x"BC8D",
    x"B07F",
    x"A57E",
    x"9BB1",
    x"9338",
    x"8C30",
    x"86B0",
    x"82CD",
    x"8092",
    x"8008",
    x"8130",
    x"8406",
    x"8881",
    x"8E92",
    x"9623",
    x"9F1C",
    x"A95D",
    x"B4C4",
    x"C12B",
    x"CE66",
    x"DC4A",
    x"EAA7",
    x"F94D",
    x"0809",
    x"16AB",
    x"24FF",
    x"32D5",
    x"4000",
    x"4C51",
    x"579F",
    x"61C3",
    x"6A9C",
    x"720C",
    x"77F8",
    x"7C4D",
    x"7EFD",
    x"7FFD",
    x"7F4B",
    x"7CEA",
    x"78E0",
    x"733D",
    x"6C12",
    x"6379",
    x"598E",
    x"4E73",
    x"424E",
    x"3548",
    x"278E",
    x"194D",
    x"0AB6",
    x"FBFB",
    x"ED4D",
    x"DEDF",
    x"D0E2",
    x"C384",
    x"B6F3",
    x"AB5B",
    x"A0E1",
    x"97AB",
    x"8FD6",
    x"897E",
    x"84B8",
    x"8194",
    x"801E",
    x"8059",
    x"8245",
    x"85DC",
    x"8B12",
    x"91D4",
    x"9A0C",
    x"A39E",
    x"AE6A",
    x"BA4A",
    x"C717",
    x"D4A5",
    x"E2C6",
    x"F14A",
    x"0000",
    x"0EB6",
    x"1D3A",
    x"2B5B",
    x"38E9",
    x"45B6",
    x"5196",
    x"5C62",
    x"65F4",
    x"6E2C",
    x"74EE",
    x"7A24",
    x"7DBB",
    x"7FA7",
    x"7FE2",
    x"7E6C",
    x"7B48",
    x"7682",
    x"702A",
    x"6855",
    x"5F1F",
    x"54A5",
    x"490D",
    x"3C7C",
    x"2F1E",
    x"2121",
    x"12B3",
    x"0405",
    x"F54A",
    x"E6B3",
    x"D872",
    x"CAB8",
    x"BDB2",
    x"B18D",
    x"A672",
    x"9C87",
    x"93EE",
    x"8CC3",
    x"8720",
    x"8316",
    x"80B5",
    x"8003",
    x"8103",
    x"83B3",
    x"8808",
    x"8DF4",
    x"9564",
    x"9E3D",
    x"A861",
    x"B3AF",
    x"C001",
    x"CD2B",
    x"DB01",
    x"E955",
    x"F7F7",
    x"06B3",
    x"1559",
    x"23B6",
    x"319A",
    x"3ED5",
    x"4B3C",
    x"56A3",
    x"60E4",
    x"69DD",
    x"716E",
    x"777F",
    x"7BFA",
    x"7ED0",
    x"7FF8",
    x"7F6E",
    x"7D33",
    x"7950",
    x"73D0",
    x"6CC8",
    x"644F",
    x"5A82",
    x"4F81",
    x"4373",
    x"3680",
    x"28D3",
    x"1A9D",
    x"0C0C",
    x"FD52",
    x"EEA1",
    x"E02B",
    x"D221",
    x"C4B3",
    x"B80E",
    x"AC5D",
    x"A1C8",
    x"9873",
    x"907D",
    x"8A01",
    x"8516",
    x"81CC",
    x"802E",
    x"8042",
    x"8207",
    x"8578",
    x"8A88",
    x"9127",
    x"993E",
    x"A2B2",
    x"AD62",
    x"B92B",
    x"C5E4",
    x"D362",
    x"E178",
    x"EFF5",
    x"FEA9",
    x"0D61",
    x"1BEC",
    x"2A18",
    x"37B5",
    x"4495",
    x"508D",
    x"5B73",
    x"6523",
    x"6D7C",
    x"7461",
    x"79BB",
    x"7D79",
    x"7F8C",
    x"7FEF",
    x"7E9F",
    x"7BA2",
    x"7702",
    x"70CE",
    x"691B",
    x"6003",
    x"55A5",
    x"4A25",
    x"3DAA",
    x"305D",
    x"226C",
    x"1406",
    x"055C",
    x"F6A0",
    x"E804",
    x"D9B9",
    x"CBF0",
    x"BED8",
    x"B29D",
    x"A769",
    x"9D61",
    x"94A7",
    x"8D5A",
    x"8792",
    x"8363",
    x"80DA",
    x"8001",
    x"80DA",
    x"8363",
    x"8792",
    x"8D5A",
    x"94A7",
    x"9D61",
    x"A769",
    x"B29D",
    x"BED8",
    x"CBF0",
    x"D9B9",
    x"E804",
    x"F6A0",
    x"055C",
    x"1406",
    x"226C",
    x"305D",
    x"3DAA",
    x"4A25",
    x"55A5",
    x"6003",
    x"691B",
    x"70CE",
    x"7702",
    x"7BA2",
    x"7E9F",
    x"7FEF",
    x"7F8C",
    x"7D79",
    x"79BB",
    x"7461",
    x"6D7C",
    x"6523",
    x"5B73",
    x"508D",
    x"4495",
    x"37B5",
    x"2A18",
    x"1BEC",
    x"0D61",
    x"FEA9",
    x"EFF5",
    x"E178",
    x"D362",
    x"C5E4",
    x"B92B",
    x"AD62",
    x"A2B2",
    x"993E",
    x"9127",
    x"8A88",
    x"8578",
    x"8207",
    x"8042",
    x"802E",
    x"81CC",
    x"8516",
    x"8A01",
    x"907D",
    x"9873",
    x"A1C8",
    x"AC5D",
    x"B80E",
    x"C4B3",
    x"D221",
    x"E02B",
    x"EEA1",
    x"FD52",
    x"0C0C",
    x"1A9D",
    x"28D3",
    x"3680",
    x"4373",
    x"4F81",
    x"5A82",
    x"644F",
    x"6CC8",
    x"73D0",
    x"7950",
    x"7D33",
    x"7F6E",
    x"7FF8",
    x"7ED0",
    x"7BFA",
    x"777F",
    x"716E",
    x"69DD",
    x"60E4",
    x"56A3",
    x"4B3C",
    x"3ED5",
    x"319A",
    x"23B6",
    x"1559",
    x"06B3",
    x"F7F7",
    x"E955",
    x"DB01",
    x"CD2B",
    x"C000",
    x"B3AF",
    x"A861",
    x"9E3D",
    x"9564",
    x"8DF4",
    x"8808",
    x"83B3",
    x"8103",
    x"8003",
    x"80B5",
    x"8316",
    x"8720",
    x"8CC3",
    x"93EE",
    x"9C87",
    x"A672",
    x"B18D",
    x"BDB2",
    x"CAB8",
    x"D872",
    x"E6B3",
    x"F54A",
    x"0405",
    x"12B3",
    x"2121",
    x"2F1E",
    x"3C7C",
    x"490D",
    x"54A5",
    x"5F1F",
    x"6855",
    x"702A",
    x"7682",
    x"7B48",
    x"7E6C",
    x"7FE2",
    x"7FA7",
    x"7DBB",
    x"7A24",
    x"74EE",
    x"6E2C",
    x"65F4",
    x"5C62",
    x"5196",
    x"45B6",
    x"38E9",
    x"2B5B",
    x"1D3A",
    x"0EB6",
    x"0000",
    x"F14A",
    x"E2C6",
    x"D4A5",
    x"C717",
    x"BA4A",
    x"AE6A",
    x"A39E",
    x"9A0C",
    x"91D4",
    x"8B12",
    x"85DC",
    x"8245",
    x"8059",
    x"801E",
    x"8194",
    x"84B8",
    x"897E",
    x"8FD6",
    x"97AB",
    x"A0E1",
    x"AB5B",
    x"B6F3",
    x"C384",
    x"D0E2",
    x"DEDF",
    x"ED4D",
    x"FBFB",
    x"0AB6",
    x"194D",
    x"278E",
    x"3548",
    x"424E",
    x"4E73",
    x"598E",
    x"6379",
    x"6C12",
    x"733D",
    x"78E0",
    x"7CEA",
    x"7F4B",
    x"7FFD",
    x"7EFD",
    x"7C4D",
    x"77F8",
    x"720C",
    x"6A9C",
    x"61C3",
    x"579F",
    x"4C51",
    x"3FFF",
    x"32D5",
    x"24FF",
    x"16AB",
    x"0809",
    x"F94D",
    x"EAA7",
    x"DC4A",
    x"CE66",
    x"C12B",
    x"B4C4",
    x"A95D",
    x"9F1C",
    x"9623",
    x"8E92",
    x"8881",
    x"8406",
    x"8130",
    x"8008",
    x"8092",
    x"82CD",
    x"86B0",
    x"8C30",
    x"9338",
    x"9BB1",
    x"A57E",
    x"B07F",
    x"BC8D",
    x"C980",
    x"D72D",
    x"E563",
    x"F3F4",
    x"02AE",
    x"115F",
    x"1FD5",
    x"2DDF",
    x"3B4D",
    x"47F2",
    x"53A3",
    x"5E38",
    x"678D",
    x"6F83",
    x"75FF",
    x"7AEA",
    x"7E34",
    x"7FD2",
    x"7FBE",
    x"7DF9",
    x"7A88",
    x"7578",
    x"6ED9",
    x"66C2",
    x"5D4E",
    x"529E",
    x"46D5",
    x"3A1C",
    x"2C9E",
    x"1E88",
    x"100B",
    x"0157",
    x"F29F",
    x"E414",
    x"D5E8",
    x"C84B",
    x"BB6B",
    x"AF73",
    x"A48D",
    x"9ADD",
    x"9284",
    x"8B9F",
    x"8645",
    x"8287",
    x"8074",
    x"8011",
    -- nota 10
    x"0000",
    x"0F95",
    x"1EEF",
    x"2DD2",
    x"3C08",
    x"4959",
    x"5592",
    x"6086",
    x"6A0A",
    x"71FA",
    x"7838",
    x"7CAC",
    x"7F46",
    x"7FFB",
    x"7EC9",
    x"7BB3",
    x"76C7",
    x"7016",
    x"67BB",
    x"5DD5",
    x"5289",
    x"4603",
    x"3872",
    x"2A0A",
    x"1B03",
    x"0B94",
    x"FBF9",
    x"EC6E",
    x"DD2D",
    x"CE71",
    x"C072",
    x"B364",
    x"A77A",
    x"9CE2",
    x"93C3",
    x"8C40",
    x"8675",
    x"827A",
    x"805D",
    x"8025",
    x"81D5",
    x"8565",
    x"8AC8",
    x"91E9",
    x"9AAE",
    x"A4F4",
    x"B095",
    x"BD65",
    x"CB32",
    x"D9C8",
    x"E8F0",
    x"F870",
    x"080C",
    x"178A",
    x"26AE",
    x"353F",
    x"4305",
    x"4FCC",
    x"5B63",
    x"659E",
    x"6E56",
    x"756A",
    x"7ABE",
    x"7E40",
    x"7FE0",
    x"7F9A",
    x"7D6D",
    x"7963",
    x"738B",
    x"6BFB",
    x"62CF",
    x"582C",
    x"4C38",
    x"3F23",
    x"311C",
    x"225B",
    x"1317",
    x"038A",
    x"F3F0",
    x"E484",
    x"D580",
    x"C71F",
    x"B995",
    x"AD18",
    x"A1D7",
    x"97FC",
    x"8FAE",
    x"890B",
    x"842D",
    x"8127",
    x"8003",
    x"80C7",
    x"8370",
    x"87F3",
    x"8E3F",
    x"963C",
    x"9FCC",
    x"AACB",
    x"B70D",
    x"C466",
    x"D2A2",
    x"E18A",
    x"F0E6",
    x"007C",
    x"1010",
    x"1F67",
    x"2E46",
    x"3C75",
    x"49BE",
    x"55EE",
    x"60D7",
    x"6A4F",
    x"7232",
    x"7862",
    x"7CC8",
    x"7F53",
    x"7FF9",
    x"7EB7",
    x"7B93",
    x"7699",
    x"6FDA",
    x"6772",
    x"5D80",
    x"522A",
    x"459B",
    x"3802",
    x"2995",
    x"1A89",
    x"0B18",
    x"FB7D",
    x"EBF3",
    x"DCB6",
    x"CDFF",
    x"C006",
    x"B301",
    x"A721",
    x"9C93",
    x"9381",
    x"8C0B",
    x"864F",
    x"8262",
    x"8054",
    x"802C",
    x"81EA",
    x"8589",
    x"8AFA",
    x"9229",
    x"9AFA",
    x"A54C",
    x"B0F7",
    x"BDCF",
    x"CBA3",
    x"DA3F",
    x"E96A",
    x"F8EC",
    x"0888",
    x"1804",
    x"2724",
    x"35B0",
    x"436F",
    x"502D",
    x"5BBA",
    x"65E9",
    x"6E95",
    x"759B",
    x"7AE1",
    x"7E54",
    x"7FE5",
    x"7F90",
    x"7D54",
    x"793C",
    x"7355",
    x"6BB8",
    x"6280",
    x"57D2",
    x"4BD4",
    x"3EB6",
    x"30AA",
    x"21E3",
    x"129C",
    x"030E",
    x"F375",
    x"E40B",
    x"D50B",
    x"C6AF",
    x"B92E",
    x"ACBA",
    x"A183",
    x"97B4",
    x"8F72",
    x"88DD",
    x"840E",
    x"8116",
    x"8002",
    x"80D5",
    x"838D",
    x"881E",
    x"8E78",
    x"9682",
    x"A01E",
    x"AB27",
    x"B774",
    x"C4D4",
    x"D316",
    x"E203",
    x"F162",
    x"00F8",
    x"108B",
    x"1FDF",
    x"2EBA",
    x"3CE3",
    x"4A24",
    x"564A",
    x"6128",
    x"6A94",
    x"726A",
    x"788C",
    x"7CE4",
    x"7F5F",
    x"7FF6",
    x"7EA5",
    x"7B73",
    x"766A",
    x"6F9E",
    x"6729",
    x"5D2B",
    x"51CA",
    x"4532",
    x"3793",
    x"291F",
    x"1A10",
    x"0A9D",
    x"FB01",
    x"EB79",
    x"DC3E",
    x"CD8C",
    x"BF9A",
    x"B29E",
    x"A6C8",
    x"9C45",
    x"933F",
    x"8BD6",
    x"8628",
    x"824A",
    x"804B",
    x"8032",
    x"8200",
    x"85AD",
    x"8B2D",
    x"9269",
    x"9B47",
    x"A5A4",
    x"B159",
    x"BE3A",
    x"CC15",
    x"DAB6",
    x"E9E5",
    x"F968",
    x"0904",
    x"187E",
    x"279B",
    x"3620",
    x"43D8",
    x"508D",
    x"5C10",
    x"6634",
    x"6ED3",
    x"75CC",
    x"7B04",
    x"7E68",
    x"7FEA",
    x"7F85",
    x"7D3B",
    x"7914",
    x"731F",
    x"6B75",
    x"6231",
    x"5777",
    x"4B70",
    x"3E4A",
    x"3037",
    x"216C",
    x"1221",
    x"0292",
    x"F2F9",
    x"E392",
    x"D496",
    x"C640",
    x"B8C7",
    x"AC5C",
    x"A130",
    x"976C",
    x"8F38",
    x"88B0",
    x"83EF",
    x"8106",
    x"8001",
    x"80E4",
    x"83AA",
    x"884A",
    x"8EB2",
    x"96C9",
    x"A071",
    x"AB85",
    x"B7DA",
    x"C542",
    x"D38A",
    x"E27B",
    x"F1DD",
    x"0175",
    x"1107",
    x"2058",
    x"2F2E",
    x"3D50",
    x"4A89",
    x"56A6",
    x"6179",
    x"6AD9",
    x"72A2",
    x"78B6",
    x"7CFF",
    x"7F6B",
    x"7FF3",
    x"7E93",
    x"7B52",
    x"763A",
    x"6F61",
    x"66DF",
    x"5CD6",
    x"516B",
    x"44CA",
    x"3723",
    x"28AA",
    x"1996",
    x"0A21",
    x"FA85",
    x"EAFE",
    x"DBC7",
    x"CD1A",
    x"BF2F",
    x"B23B",
    x"A66F",
    x"9BF8",
    x"92FE",
    x"8BA2",
    x"8603",
    x"8233",
    x"8043",
    x"8039",
    x"8216",
    x"85D2",
    x"8B60",
    x"92A9",
    x"9B93",
    x"A5FC",
    x"B1BB",
    x"BEA4",
    x"CC86",
    x"DB2D",
    x"EA5F",
    x"F9E4",
    x"0980",
    x"18F8",
    x"2811",
    x"3691",
    x"4441",
    x"50EE",
    x"5C66",
    x"667F",
    x"6F11",
    x"75FC",
    x"7B26",
    x"7E7B",
    x"7FEE",
    x"7F7A",
    x"7D21",
    x"78EB",
    x"72E9",
    x"6B31",
    x"61E1",
    x"571C",
    x"4B0C",
    x"3DDD",
    x"2FC3",
    x"20F4",
    x"11A6",
    x"0216",
    x"F27D",
    x"E319",
    x"D422",
    x"C5D2",
    x"B85F",
    x"ABFE",
    x"A0DC",
    x"9725",
    x"8EFD",
    x"8883",
    x"83D1",
    x"80F7",
    x"8001",
    x"80F2",
    x"83C8",
    x"8876",
    x"8EEC",
    x"9710",
    x"A0C4",
    x"ABE2",
    x"B841",
    x"C5B1",
    x"D3FF",
    x"E2F4",
    x"F259",
    x"01F1",
    x"1182",
    x"20D0",
    x"2FA1",
    x"3DBD",
    x"4AEE",
    x"5701",
    x"61C9",
    x"6B1D",
    x"72D9",
    x"78DF",
    x"7D19",
    x"7F77",
    x"7FEF",
    x"7E81",
    x"7B30",
    x"760A",
    x"6F23",
    x"6695",
    x"5C80",
    x"510B",
    x"4461",
    x"36B2",
    x"2834",
    x"191C",
    x"09A5",
    x"FA09",
    x"EA84",
    x"DB50",
    x"CCA8",
    x"BEC4",
    x"B1D8",
    x"A616",
    x"9BAA",
    x"92BD",
    x"8B6F",
    x"85DD",
    x"821D",
    x"803B",
    x"8041",
    x"822C",
    x"85F7",
    x"8B93",
    x"92EA",
    x"9BE1",
    x"A654",
    x"B21D",
    x"BF0F",
    x"CCF8",
    x"DBA4",
    x"EADA",
    x"FA60",
    x"09FC",
    x"1972",
    x"2887",
    x"3701",
    x"44AA",
    x"514E",
    x"5CBC",
    x"66C9",
    x"6F4E",
    x"762C",
    x"7B48",
    x"7E8E",
    x"7FF2",
    x"7F6F",
    x"7D07",
    x"78C2",
    x"72B2",
    x"6AED",
    x"6191",
    x"56C1",
    x"4AA7",
    x"3D70",
    x"2F50",
    x"207C",
    x"112B",
    x"019A",
    x"F202",
    x"E2A0",
    x"D3AD",
    x"C563",
    x"B7F9",
    x"ABA0",
    x"A089",
    x"96DE",
    x"8EC3",
    x"8857",
    x"83B3",
    x"80E8",
    x"8001",
    x"8102",
    x"83E6",
    x"88A3",
    x"8F26",
    x"9757",
    x"A117",
    x"AC40",
    x"B8A8",
    x"C61F",
    x"D474",
    x"E36D",
    x"F2D4",
    x"026D",
    x"11FD",
    x"2148",
    x"3014",
    x"3E2A",
    x"4B52",
    x"575C",
    x"6219",
    x"6B61",
    x"730F",
    x"7908",
    x"7D33",
    x"7F82",
    x"7FEB",
    x"7E6D",
    x"7B0E",
    x"75DA",
    x"6EE5",
    x"664A",
    x"5C2A",
    x"50AA",
    x"43F8",
    x"3642",
    x"27BE",
    x"18A2",
    x"0929",
    x"F98D",
    x"EA09",
    x"DAD9",
    x"CC37",
    x"BE59",
    x"B176",
    x"A5BE",
    x"9B5D",
    x"927C",
    x"8B3C",
    x"85B8",
    x"8206",
    x"8034",
    x"8049",
    x"8243",
    x"861D",
    x"8BC7",
    x"932B",
    x"9C2E",
    x"A6AD",
    x"B280",
    x"BF7A",
    x"CD6A",
    x"DC1B",
    x"EB54",
    x"FADC",
    x"0A78",
    x"19EB",
    x"28FC",
    x"3771",
    x"4513",
    x"51AE",
    x"5D11",
    x"6713",
    x"6F8B",
    x"765B",
    x"7B69",
    x"7EA0",
    x"7FF5",
    x"7F63",
    x"7CEC",
    x"7899",
    x"727B",
    x"6AA8",
    x"6140",
    x"5665",
    x"4A42",
    x"3D03",
    x"2EDD",
    x"2003",
    x"10B0",
    x"011D",
    x"F187",
    x"E227",
    x"D339",
    x"C4F5",
    x"B792",
    x"AB43",
    x"A037",
    x"9697",
    x"8E89",
    x"882B",
    x"8395",
    x"80DA",
    x"8002",
    x"8111",
    x"8405",
    x"88D0",
    x"8F61",
    x"979F",
    x"A16A",
    x"AC9E",
    x"B90F",
    x"C68E",
    x"D4E8",
    x"E3E7",
    x"F350",
    x"02E9",
    x"1278",
    x"21C0",
    x"3087",
    x"3E96",
    x"4BB6",
    x"57B7",
    x"6269",
    x"6BA4",
    x"7345",
    x"7930",
    x"7D4D",
    x"7F8D",
    x"7FE7",
    x"7E5A",
    x"7AEC",
    x"75A9",
    x"6EA7",
    x"6600",
    x"5BD3",
    x"504A",
    x"438E",
    x"35D1",
    x"2748",
    x"1828",
    x"08AD",
    x"F911",
    x"E98F",
    x"DA62",
    x"CBC5",
    x"BDEF",
    x"B114",
    x"A566",
    x"9B11",
    x"923C",
    x"8B09",
    x"8594",
    x"81F1",
    x"802D",
    x"8051",
    x"825B",
    x"8643",
    x"8BFB",
    x"936D",
    x"9C7C",
    x"A706",
    x"B2E3",
    x"BFE6",
    x"CDDC",
    x"DC92",
    x"EBCF",
    x"FB58",
    x"0AF3",
    x"1A65",
    x"2972",
    x"37E1",
    x"457B",
    x"520D",
    x"5D67",
    x"675C",
    x"6FC8",
    x"768B",
    x"7B89",
    x"7EB2",
    x"7FF8",
    x"7F57",
    x"7CD1",
    x"786F",
    x"7243",
    x"6A64",
    x"60EF",
    x"560A",
    x"49DD",
    x"3C96",
    x"2E69",
    x"1F8B",
    x"1035",
    x"00A1",
    x"F10B",
    x"E1AE",
    x"D2C4",
    x"C487",
    x"B72C",
    x"AAE6",
    x"9FE5",
    x"9651",
    x"8E50",
    x"8800",
    x"8378",
    x"80CC",
    x"8003",
    x"8122",
    x"8424",
    x"88FD",
    x"8F9C",
    x"97E7",
    x"A1BE",
    x"ACFC",
    x"B977",
    x"C6FD",
    x"D55D",
    x"E460",
    x"F3CB",
    x"0365",
    x"12F3",
    x"2237",
    x"30FA",
    x"3F02",
    x"4C1A",
    x"5811",
    x"62B8",
    x"6BE7",
    x"737B",
    x"7958",
    x"7D66",
    x"7F97",
    x"7FE2",
    x"7E46",
    x"7AC9",
    x"7578",
    x"6E69",
    x"65B4",
    x"5B7D",
    x"4FE9",
    x"4325",
    x"3561",
    x"26D1",
    x"17AE",
    x"0831",
    x"F895",
    x"E915",
    x"D9EC",
    x"CB54",
    x"BD85",
    x"B0B3",
    x"A50E",
    x"9AC5",
    x"91FC",
    x"8AD7",
    x"8570",
    x"81DB",
    x"8027",
    x"805A",
    x"8273",
    x"866A",
    x"8C30",
    x"93AF",
    x"9CCA",
    x"A760",
    x"B346",
    x"C051",
    x"CE4F",
    x"DD0A",
    x"EC49",
    x"FBD4",
    x"0B6F",
    x"1ADE",
    x"29E7",
    x"3851",
    x"45E4",
    x"526C",
    x"5DBB",
    x"67A5",
    x"7005",
    x"76B9",
    x"7BAA",
    x"7EC3",
    x"7FFA",
    x"7F4A",
    x"7CB5",
    x"7845",
    x"720B",
    x"6A1E",
    x"609E",
    x"55AE",
    x"4977",
    x"3C29",
    x"2DF5",
    x"1F13",
    x"0FBA",
    x"0025",
    x"F090",
    x"E135",
    x"D250",
    x"C419",
    x"B6C6",
    x"AA8A",
    x"9F93",
    x"960B",
    x"8E17",
    x"87D5",
    x"835C",
    x"80BE",
    x"8004",
    x"8132",
    x"8443",
    x"892B",
    x"8FD8",
    x"982F",
    x"A212",
    x"AD5B",
    x"B9DE",
    x"C76D",
    x"D5D3",
    x"E4D9",
    x"F447",
    x"03E2",
    x"136D",
    x"22AF",
    x"316D",
    x"3F6E",
    x"4C7E",
    x"586B",
    x"6307",
    x"6C2A",
    x"73B1",
    x"797F",
    x"7D7F",
    x"7FA0",
    x"7FDC",
    x"7E31",
    x"7AA5",
    x"7547",
    x"6E29",
    x"6569",
    x"5B26",
    x"4F88",
    x"42BB",
    x"34F0",
    x"265B",
    x"1734",
    x"07B5",
    x"F819",
    x"E89A",
    x"D975",
    x"CAE3",
    x"BD1B",
    x"B051",
    x"A4B7",
    x"9A79",
    x"91BD",
    x"8AA5",
    x"854C",
    x"81C7",
    x"8021",
    x"8063",
    x"828B",
    x"8691",
    x"8C65",
    x"93F1",
    x"9D19",
    x"A7B9",
    x"B3AA",
    x"C0BD",
    x"CEC1",
    x"DD81",
    x"ECC4",
    x"FC51",
    x"0BEB",
    x"1B58",
    x"2A5D",
    x"38C0",
    x"464C",
    x"52CB",
    x"5E10",
    x"67EE",
    x"7040",
    x"76E7",
    x"7BCA",
    x"7ED4",
    x"7FFC",
    x"7F3D",
    x"7C99",
    x"781A",
    x"71D2",
    x"69D9",
    x"604C",
    x"5551",
    x"4911",
    x"3BBB",
    x"2D81",
    x"1E9A",
    x"0F3E",
    x"FFA9",
    x"F015",
    x"E0BD",
    x"D1DC",
    x"C3AB",
    x"B660",
    x"AA2D",
    x"9F41",
    x"95C6",
    x"8DDF",
    x"87AA",
    x"8340",
    x"80B1",
    x"8007",
    x"8144",
    x"8463",
    x"895A",
    x"9014",
    x"9878",
    x"A267",
    x"ADBA",
    x"BA46",
    x"C7DC",
    x"D648",
    x"E553",
    x"F4C3",
    x"045E",
    x"13E8",
    x"2327",
    x"31DF",
    x"3FDA",
    x"4CE2",
    x"58C4",
    x"6355",
    x"6C6C",
    x"73E5",
    x"79A6",
    x"7D97",
    x"7FAA",
    x"7FD6",
    x"7E1C",
    x"7A82",
    x"7515",
    x"6DEA",
    x"651D",
    x"5ACE",
    x"4F26",
    x"4251",
    x"347E",
    x"25E4",
    x"16BA",
    x"0739",
    x"F79D",
    x"E820",
    x"D8FF",
    x"CA72",
    x"BCB1",
    x"AFF0",
    x"A460",
    x"9A2D",
    x"917E",
    x"8A74",
    x"8529",
    x"81B2",
    x"801C",
    x"806D",
    x"82A4",
    x"86B8",
    x"8C9A",
    x"9434",
    x"9D68",
    x"A814",
    x"B40E",
    x"C129",
    x"CF34",
    x"DDF9",
    x"ED3F",
    x"FCCD",
    x"0C67",
    x"1BD1",
    x"2AD2",
    x"392F",
    x"46B3",
    x"532A",
    x"5E64",
    x"6836",
    x"707C",
    x"7715",
    x"7BE9",
    x"7EE5",
    x"7FFE",
    x"7F2F",
    x"7C7C",
    x"77EF",
    x"7199",
    x"6993",
    x"5FFA",
    x"54F4",
    x"48AB",
    x"3B4D",
    x"2D0D",
    x"1E21",
    x"0EC3",
    x"FF2D",
    x"EF99",
    x"E044",
    x"D168",
    x"C33E",
    x"B5FB",
    x"A9D1",
    x"9EF0",
    x"9581",
    x"8DA7",
    x"8780",
    x"8324",
    x"80A4",
    x"8009",
    x"8155",
    x"8484",
    x"8988",
    x"9050",
    x"98C1",
    x"A2BC",
    -- nota 11
    x"0000",
    x"1081",
    x"20BB",
    x"306A",
    x"3F49",
    x"4D1A",
    x"59A2",
    x"64AA",
    x"6E05",
    x"7589",
    x"7B17",
    x"7E96",
    x"7FF9",
    x"7F39",
    x"7C59",
    x"7765",
    x"7074",
    x"67A1",
    x"5D14",
    x"50F9",
    x"4384",
    x"34EF",
    x"2577",
    x"155F",
    x"04EC",
    x"F463",
    x"E40D",
    x"D42E",
    x"C50A",
    x"B6E2",
    x"A9F2",
    x"9E73",
    x"9494",
    x"8C80",
    x"865A",
    x"823C",
    x"8037",
    x"8055",
    x"8294",
    x"86EB",
    x"8D48",
    x"958F",
    x"9F9D",
    x"AB46",
    x"B85A",
    x"C6A0",
    x"D5DC",
    x"E5CB",
    x"F62A",
    x"06B4",
    x"1721",
    x"272B",
    x"368D",
    x"4507",
    x"5259",
    x"5E4B",
    x"68AB",
    x"714B",
    x"7807",
    x"7CC2",
    x"7F68",
    x"7FED",
    x"7E50",
    x"7A96",
    x"74D1",
    x"6D19",
    x"638E",
    x"585A",
    x"4BAC",
    x"3DBB",
    x"2EC2",
    x"1F01",
    x"0EBC",
    x"FE37",
    x"EDBB",
    x"DD8C",
    x"CDF1",
    x"BF2B",
    x"B17B",
    x"A51A",
    x"9A3E",
    x"9115",
    x"89C5",
    x"846F",
    x"8129",
    x"8001",
    x"80FD",
    x"8417",
    x"8942",
    x"9069",
    x"996D",
    x"A428",
    x"B06A",
    x"BE01",
    x"CCB2",
    x"DC3F",
    x"EC64",
    x"FCDD",
    x"0D63",
    x"1DB0",
    x"2D7E",
    x"3C8A",
    x"4A93",
    x"575E",
    x"62B3",
    x"6C62",
    x"7442",
    x"7A31",
    x"7E16",
    x"7FE0",
    x"7F87",
    x"7D0E",
    x"787E",
    x"71EB",
    x"6971",
    x"5F34",
    x"5361",
    x"4629",
    x"37C6",
    x"2874",
    x"1875",
    x"080E",
    x"F784",
    x"E71F",
    x"D724",
    x"C7D7",
    x"B97B",
    x"AC4B",
    x"A082",
    x"9651",
    x"8DE3",
    x"875D",
    x"82DB",
    x"8070",
    x"8025",
    x"81FD",
    x"85F0",
    x"8BED",
    x"93D9",
    x"9D94",
    x"A8F3",
    x"B5C6",
    x"C3D7",
    x"D2E9",
    x"E2BB",
    x"F30A",
    x"0391",
    x"1409",
    x"242B",
    x"33B2",
    x"425D",
    x"4FEC",
    x"5C25",
    x"66D5",
    x"6FCD",
    x"76E7",
    x"7C05",
    x"7F11",
    x"7FFE",
    x"7EC8",
    x"7B74",
    x"7610",
    x"6EB4",
    x"657F",
    x"5A98",
    x"4E2E",
    x"4076",
    x"31AA",
    x"220A",
    x"11D8",
    x"015B",
    x"F0D7",
    x"E094",
    x"D0D8",
    x"C1E5",
    x"B3FB",
    x"A757",
    x"9C2D",
    x"92AE",
    x"8B02",
    x"854A",
    x"819F",
    x"8010",
    x"80A3",
    x"8357",
    x"881F",
    x"8EE8",
    x"9795",
    x"A1FF",
    x"ADFB",
    x"BB56",
    x"C9D7",
    x"D93E",
    x"E94C",
    x"F9BA",
    x"0A43",
    x"1AA1",
    x"2A8C",
    x"39C2",
    x"4801",
    x"550C",
    x"60AC",
    x"6AAE",
    x"72E9",
    x"7938",
    x"7D82",
    x"7FB3",
    x"7FC2",
    x"7DAF",
    x"7983",
    x"7350",
    x"6B30",
    x"6146",
    x"55BC",
    x"48C4",
    x"3A95",
    x"2B6B",
    x"1B88",
    x"0B2F",
    x"FAA6",
    x"EA34",
    x"DA20",
    x"CAAD",
    x"BC1E",
    x"AEB2",
    x"A2A0",
    x"981E",
    x"8F58",
    x"8873",
    x"838D",
    x"80BB",
    x"8009",
    x"817A",
    x"8508",
    x"8AA3",
    x"9234",
    x"9B9A",
    x"A6AD",
    x"B33E",
    x"C117",
    x"CFFC",
    x"DFAF",
    x"EFEC",
    x"006E",
    x"10EE",
    x"2126",
    x"30D0",
    x"3FA9",
    x"4D72",
    x"59F0",
    x"64EE",
    x"6E3D",
    x"75B4",
    x"7B35",
    x"7EA6",
    x"7FFB",
    x"7F2C",
    x"7C3E",
    x"773D",
    x"703F",
    x"6761",
    x"5CC9",
    x"50A4",
    x"4327",
    x"348A",
    x"250D",
    x"14F2",
    x"047E",
    x"F3F6",
    x"E3A1",
    x"D3C6",
    x"C4A8",
    x"B687",
    x"A9A1",
    x"9E2B",
    x"9458",
    x"8C51",
    x"8638",
    x"8228",
    x"8031",
    x"805D",
    x"82AA",
    x"870F",
    x"8D79",
    x"95CC",
    x"9FE5",
    x"AB99",
    x"B8B6",
    x"C703",
    x"D644",
    x"E637",
    x"F698",
    x"0722",
    x"178D",
    x"2793",
    x"36F1",
    x"4563",
    x"52AD",
    x"5E96",
    x"68EA",
    x"717E",
    x"782D",
    x"7CDA",
    x"7F72",
    x"7FE9",
    x"7E3E",
    x"7A76",
    x"74A4",
    x"6CDF",
    x"6349",
    x"580A",
    x"4B53",
    x"3D5A",
    x"2E5B",
    x"1E96",
    x"0E4E",
    x"FDC9",
    x"ED4E",
    x"DD22",
    x"CD8B",
    x"BECC",
    x"B124",
    x"A4CD",
    x"99FB",
    x"90DE",
    x"899B",
    x"8453",
    x"811B",
    x"8001",
    x"810A",
    x"8432",
    x"896B",
    x"909F",
    x"99AF",
    x"A474",
    x"B0C1",
    x"BE60",
    x"CD17",
    x"DCA9",
    x"ECD1",
    x"FD4B",
    x"0DD1",
    x"1E1B",
    x"2DE5",
    x"3CEB",
    x"4AED",
    x"57AE",
    x"62F9",
    x"6C9C",
    x"7470",
    x"7A51",
    x"7E28",
    x"7FE4",
    x"7F7E",
    x"7CF6",
    x"7858",
    x"71B8",
    x"6932",
    x"5EEB",
    x"530D",
    x"45CD",
    x"3763",
    x"280B",
    x"1809",
    x"07A0",
    x"F716",
    x"E6B3",
    x"D6BB",
    x"C774",
    x"B91F",
    x"ABF8",
    x"A039",
    x"9613",
    x"8DB2",
    x"8739",
    x"82C4",
    x"8067",
    x"802B",
    x"8211",
    x"8611",
    x"8C1B",
    x"9414",
    x"9DDA",
    x"A944",
    x"B620",
    x"C438",
    x"D350",
    x"E326",
    x"F378",
    x"03FF",
    x"1476",
    x"2495",
    x"3417",
    x"42BB",
    x"5042",
    x"5C71",
    x"6716",
    x"7002",
    x"770F",
    x"7C20",
    x"7F1E",
    x"7FFD",
    x"7EB8",
    x"7B57",
    x"75E6",
    x"6E7D",
    x"653C",
    x"5A4A",
    x"4DD7",
    x"4016",
    x"3144",
    x"21A0",
    x"116B",
    x"00EC",
    x"F06A",
    x"E02A",
    x"D071",
    x"C185",
    x"B3A3",
    x"A707",
    x"9BE8",
    x"9275",
    x"8AD6",
    x"852B",
    x"818E",
    x"800C",
    x"80AE",
    x"8370",
    x"8846",
    x"8F1C",
    x"97D5",
    x"A24A",
    x"AE50",
    x"BBB3",
    x"CA3A",
    x"D9A7",
    x"E9B8",
    x"FA28",
    x"0AB1",
    x"1B0C",
    x"2AF4",
    x"3A24",
    x"485C",
    x"555E",
    x"60F4",
    x"6AEB",
    x"7319",
    x"795B",
    x"7D97",
    x"7FBA",
    x"7FBB",
    x"7D9A",
    x"7961",
    x"7320",
    x"6AF4",
    x"60FE",
    x"556A",
    x"4869",
    x"3A33",
    x"2B03",
    x"1B1C",
    x"0AC1",
    x"FA38",
    x"E9C8",
    x"D9B7",
    x"CA49",
    x"BBC1",
    x"AE5D",
    x"A255",
    x"97DE",
    x"8F24",
    x"884C",
    x"8374",
    x"80B0",
    x"800C",
    x"818B",
    x"8527",
    x"8ACF",
    x"926C",
    x"9BDE",
    x"A6FC",
    x"B396",
    x"C177",
    x"D062",
    x"E01A",
    x"F05A",
    x"00DC",
    x"115B",
    x"2190",
    x"3135",
    x"4008",
    x"4DCA",
    x"5A3F",
    x"6532",
    x"6E75",
    x"75DF",
    x"7B52",
    x"7EB6",
    x"7FFC",
    x"7F20",
    x"7C24",
    x"7715",
    x"700A",
    x"6720",
    x"5C7D",
    x"504E",
    x"42C9",
    x"3426",
    x"24A4",
    x"1486",
    x"0410",
    x"F388",
    x"E336",
    x"D35F",
    x"C446",
    x"B62D",
    x"A950",
    x"9DE5",
    x"941D",
    x"8C22",
    x"8616",
    x"8214",
    x"802C",
    x"8065",
    x"82C1",
    x"8733",
    x"8DAA",
    x"960A",
    x"A02E",
    x"ABEC",
    x"B911",
    x"C766",
    x"D6AC",
    x"E6A3",
    x"F706",
    x"0790",
    x"17F9",
    x"27FC",
    x"3754",
    x"45C0",
    x"5301",
    x"5EE0",
    x"6929",
    x"71B1",
    x"7853",
    x"7CF2",
    x"7F7C",
    x"7FE5",
    x"7E2B",
    x"7A56",
    x"7476",
    x"6CA5",
    x"6303",
    x"57BA",
    x"4AFA",
    x"3CF9",
    x"2DF4",
    x"1E2B",
    x"0DE1",
    x"FD5B",
    x"ECE1",
    x"DCB8",
    x"CD26",
    x"BE6E",
    x"B0CD",
    x"A480",
    x"99B9",
    x"90A7",
    x"8972",
    x"8437",
    x"810C",
    x"8001",
    x"8119",
    x"844F",
    x"8995",
    x"90D6",
    x"99F2",
    x"A4C2",
    x"B117",
    x"BEBF",
    x"CD7D",
    x"DD12",
    x"ED3E",
    x"FDB9",
    x"0E3E",
    x"1E86",
    x"2E4C",
    x"3D4C",
    x"4B46",
    x"57FE",
    x"633E",
    x"6CD6",
    x"749D",
    x"7A72",
    x"7E3B",
    x"7FE9",
    x"7F74",
    x"7CDE",
    x"7833",
    x"7186",
    x"68F3",
    x"5EA1",
    x"52B9",
    x"4571",
    x"36FF",
    x"27A3",
    x"179D",
    x"0732",
    x"F6A8",
    x"E647",
    x"D653",
    x"C711",
    x"B8C3",
    x"ABA5",
    x"9FF0",
    x"95D5",
    x"8D80",
    x"8714",
    x"82AE",
    x"805E",
    x"8030",
    x"8225",
    x"8633",
    x"8C4A",
    x"944F",
    x"9E21",
    x"A995",
    x"B67A",
    x"C49A",
    x"D3B7",
    x"E392",
    x"F3E6",
    x"046D",
    x"14E2",
    x"24FE",
    x"347C",
    x"4319",
    x"5097",
    x"5CBD",
    x"6757",
    x"7037",
    x"7738",
    x"7C3B",
    x"7F2B",
    x"7FFB",
    x"7EA9",
    x"7B39",
    x"75BB",
    x"6E45",
    x"64F8",
    x"59FC",
    x"4D7F",
    x"3FB7",
    x"30DF",
    x"2135",
    x"10FE",
    x"007E",
    x"EFFC",
    x"DFBF",
    x"D00B",
    x"C125",
    x"B34B",
    x"A6B8",
    x"9BA4",
    x"923C",
    x"8AA9",
    x"850C",
    x"817D",
    x"800A",
    x"80BA",
    x"838A",
    x"886D",
    x"8F50",
    x"9815",
    x"A295",
    x"AEA5",
    x"BC11",
    x"CA9E",
    x"DA10",
    x"EA25",
    x"FA96",
    x"0B1F",
    x"1B78",
    x"2B5C",
    x"3A86",
    x"48B7",
    x"55B0",
    x"613B",
    x"6B27",
    x"7349",
    x"797E",
    x"7DAC",
    x"7FC1",
    x"7FB4",
    x"7D85",
    x"793D",
    x"72F0",
    x"6AB7",
    x"60B6",
    x"5518",
    x"480E",
    x"39D0",
    x"2A9B",
    x"1AB0",
    x"0A53",
    x"F9CA",
    x"E95C",
    x"D94E",
    x"C9E5",
    x"BB64",
    x"AE08",
    x"A20A",
    x"979E",
    x"8EF0",
    x"8825",
    x"835B",
    x"80A5",
    x"800F",
    x"819C",
    x"8546",
    x"8AFC",
    x"92A6",
    x"9C23",
    x"A74B",
    x"B3EE",
    x"C1D7",
    x"D0C9",
    x"E085",
    x"F0C7",
    x"014A",
    x"11C8",
    x"21FA",
    x"319B",
    x"4068",
    x"4E21",
    x"5A8D",
    x"6575",
    x"6EAC",
    x"760A",
    x"7B70",
    x"7EC6",
    x"7FFE",
    x"7F13",
    x"7C09",
    x"76ED",
    x"6FD4",
    x"66DE",
    x"5C30",
    x"4FF8",
    x"426B",
    x"33C1",
    x"243A",
    x"1419",
    x"03A1",
    x"F31A",
    x"E2CB",
    x"D2F8",
    x"C3E5",
    x"B5D3",
    x"A8FF",
    x"9D9E",
    x"93E2",
    x"8BF3",
    x"85F5",
    x"8200",
    x"8026",
    x"806E",
    x"82D8",
    x"8758",
    x"8DDC",
    x"9648",
    x"A077",
    x"AC3F",
    x"B96D",
    x"C7C9",
    x"D714",
    x"E70F",
    x"F774",
    x"07FE",
    x"1865",
    x"2865",
    x"37B7",
    x"461C",
    x"5355",
    x"5F2A",
    x"6968",
    x"71E3",
    x"7878",
    x"7D0A",
    x"7F86",
    x"7FE0",
    x"7E18",
    x"7A36",
    x"7448",
    x"6C6A",
    x"62BD",
    x"5769",
    x"4AA0",
    x"3C98",
    x"2D8E",
    x"1DC0",
    x"0D73",
    x"FCED",
    x"EC74",
    x"DC4E",
    x"CCC1",
    x"BE0F",
    x"B077",
    x"A433",
    x"9977",
    x"9071",
    x"8948",
    x"841B",
    x"80FF",
    x"8001",
    x"8127",
    x"846B",
    x"89BF",
    x"910D",
    x"9A34",
    x"A50F",
    x"B16E",
    x"BF1D",
    x"CDE2",
    x"DD7D",
    x"EDAB",
    x"FE27",
    x"0EAC",
    x"1EF1",
    x"2EB3",
    x"3DAD",
    x"4B9F",
    x"584E",
    x"6384",
    x"6D10",
    x"74CA",
    x"7A92",
    x"7E4D",
    x"7FEC",
    x"7F69",
    x"7CC6",
    x"780D",
    x"7153",
    x"68B4",
    x"5E56",
    x"5265",
    x"4514",
    x"369C",
    x"273A",
    x"1731",
    x"06C4",
    x"F63B",
    x"E5DB",
    x"D5EB",
    x"C6AF",
    x"B868",
    x"AB53",
    x"9FA7",
    x"9598",
    x"8D4F",
    x"86F1",
    x"8297",
    x"8056",
    x"8037",
    x"8239",
    x"8655",
    x"8C79",
    x"948B",
    x"9E68",
    x"A9E6",
    x"B6D4",
    x"C4FB",
    x"D41E",
    x"E3FD",
    x"F453",
    x"04DC",
    x"154F",
    x"2567",
    x"34E0",
    x"4377",
    x"50ED",
    x"5D09",
    x"6798",
    x"706C",
    x"7760",
    x"7C55",
    x"7F37",
    x"7FF9",
    x"7E99",
    x"7B1B",
    x"758F",
    x"6E0D",
    x"64B4",
    x"59AD",
    x"4D27",
    x"3F57",
    x"3079",
    x"20CB",
    x"1091",
    x"0010",
    x"EF8F",
    x"DF54",
    x"CFA5",
    x"C0C5",
    x"B2F2",
    x"A66A",
    x"9B60",
    x"9204",
    x"8A7E",
    x"84EE",
    x"816C",
    x"8007",
    x"80C6",
    x"83A3",
    x"8895",
    x"8F85",
    x"9855",
    x"A2E1",
    x"AEFA",
    x"BC6E",
    x"CB03",
    x"DA7A",
    x"EA91",
    x"FB04",
    x"0B8D",
    x"1BE4",
    x"2BC3",
    x"3AE8",
    x"4911",
    x"5602",
    x"6183",
    x"6B63",
    x"7379",
    x"79A1",
    x"7DC1",
    x"7FC8",
    x"7FAC",
    x"7D6F",
    x"791A",
    x"72BF",
    x"6A7A",
    x"606E",
    x"54C6",
    x"47B3",
    x"396E",
    x"2A34",
    x"1A45",
    x"09E6",
    x"F95C",
    x"E8EF",
    x"D8E5",
    x"C981",
    x"BB07",
    x"ADB3",
    x"A1BF",
    x"975E",
    x"8EBC",
    x"87FF",
    x"8342",
    x"809A",
    x"8012",
    x"81AE",
    x"8565",
    x"8B28",
    x"92DF",
    x"9C68",
    x"A79B",
    x"B447",
    x"C237",
    x"D12F",
    x"E0EF",
    x"F134",
    x"01B9",
    x"1235",
    x"2264",
    x"3200",
    x"40C7",
    x"4E78",
    x"5ADA",
    x"65B8",
    x"6EE3",
    x"7635",
    x"7B8D",
    x"7ED5",
    x"7FFE",
    x"7F05",
    x"7BED",
    x"76C4",
    x"6F9F",
    x"669C",
    x"5BE4",
    x"4FA2",
    x"420C",
    x"335C",
    x"23D1",
    x"13AC",
    x"0333",
    x"F2AD",
    x"E25F",
    x"D291",
    x"C384",
    x"B57A",
    x"A8AE",
    x"9D58",
    x"93A7",
    x"8BC5",
    x"85D4",
    x"81ED",
    x"8021",
    x"8077",
    x"82EF",
    x"877D",
    x"8E0E",
    x"9686",
    x"A0C1",
    x"AC93",
    x"B9C9",
    x"C82C",
    x"D77D",
    x"E77B",
    x"F7E2",
    x"086C",
    x"18D1",
    x"28CD",
    -- nota 12
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    -- nota 13
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    -- nota 14
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    -- nota 15
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000",
    x"0000");
						 
begin
  addr <= nota & counter;
  process(clock) is
  begin
    if rising_edge(clock) then
      sample <= rom(to_integer(unsigned(addr)));
    end if;
  end process;
end v1;




